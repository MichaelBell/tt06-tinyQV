.lib '/home/mdb36/tt/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice' tt
