* NGSPICE file created from tt_um_MichaelBell_tinyQV.ext - technology: sky130A

.subckt sky130_fd_sc_hd__decap_3 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=0.59
.ends

.subckt sky130_fd_sc_hd__dfxtp_1 Q CLK D VPB VNB VPWR VGND
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X9 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X10 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X16 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X17 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X18 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X19 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X20 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X21 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X22 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X23 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_2 VPB VNB VGND VPWR B Y A
X0 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_1 VPB VNB VGND VPWR X A B
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_1 VPB VNB VGND VPWR A Y B
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2_1 VPWR VGND X B A VPB VNB
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3_1 VGND VPWR X B A C VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 VGND VPWR X A VPB VNB
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3b_1 VGND VPWR VPB VNB B C_N A X
X0 a_109_93# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 a_215_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VGND a_109_93# a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND A a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 VPWR A a_369_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 a_369_297# B a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_215_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X7 a_297_297# a_109_93# a_215_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_109_93# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 X a_215_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlygate4sd3_1 X A VPB VNB VGND VPWR
X0 VPWR A a_49_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 VGND a_285_47# a_391_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.5
X2 X a_391_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3 VGND A a_49_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VPWR a_285_47# a_391_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.5
X5 a_285_47# a_49_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X6 a_285_47# a_49_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X7 X a_391_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_1 VPWR VGND VPB VNB A2 A1 B1 Y
X0 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X3 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X4 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_6 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.97
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.05
.ends

.subckt sky130_fd_sc_hd__dlygate4sd1_1 VPWR VGND VPB VNB X A
X0 X a_299_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X1 VPWR a_193_47# a_299_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 VGND a_193_47# a_299_93# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 X a_299_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X7 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_8 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=2.89
.ends

.subckt sky130_fd_sc_hd__a21o_1 VPWR VGND VPB VNB A2 A1 B1 X
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux2_1 VGND VPWR VPB VNB X A1 S A0
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux2_2 VGND VPWR VPB VNB S A1 A0 X
X0 VPWR S a_591_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0672 ps=0.85 w=0.64 l=0.15
X1 a_591_369# A0 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1312 ps=1.05 w=0.64 l=0.15
X2 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1778 pd=1.415 as=0.135 ps=1.27 w=1 l=0.15
X3 a_79_21# A1 a_306_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1312 pd=1.05 as=0.2288 ps=1.355 w=0.64 l=0.15
X4 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND S a_578_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.05775 ps=0.695 w=0.42 l=0.15
X6 a_306_369# a_257_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2288 pd=1.355 as=0.1778 ps=1.415 w=0.64 l=0.15
X7 a_79_21# A0 a_288_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17325 pd=1.245 as=0.06825 ps=0.745 w=0.42 l=0.15
X8 a_288_47# a_257_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.097 ps=0.975 w=0.42 l=0.15
X9 a_257_199# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_578_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.17325 ps=1.245 w=0.42 l=0.15
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 a_257_199# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1728 pd=1.82 as=0.0864 ps=0.91 w=0.64 l=0.15
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__xor2_1 VNB VPB VPWR VGND A X B
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211o_1 VNB VPB VGND VPWR X A2 B1 A1 C1
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1 a_80_21# C1 a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X2 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X5 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X6 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_80_21# A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 a_472_297# B1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X9 a_80_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ai_1 VGND VPWR A2 B1 Y A1 VPB VNB
X0 Y A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X3 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_6 VPWR VGND X A VPB VNB
X0 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_161_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A a_161_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VPWR A a_161_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_161_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_4 VPB VNB VGND VPWR B Y A
X0 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3_4 VNB VPB VGND VPWR C A Y B
X0 a_27_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_27_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 Y A a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 Y A a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_27_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_27_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 a_445_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12 a_445_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VGND C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_445_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X17 a_445_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X22 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X23 VGND C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfxtp_2 Q CLK D VPB VNB VPWR VGND
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2 VPWR a_1059_315# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X4 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X8 VGND a_1059_315# Q VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X13 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X14 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X16 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X18 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X19 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X20 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X21 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X22 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X23 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X24 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X25 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 VGND VPWR A X VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211a_1 VNB VPB VGND VPWR X A1 A2 B1 C1
X0 VGND A1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_510_47# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X2 a_79_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X3 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X4 a_79_21# A2 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.1625 ps=1.325 w=1 l=0.15
X5 a_297_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X6 a_79_21# C1 a_510_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.11375 ps=1 w=0.65 l=0.15
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9 a_215_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.105625 ps=0.975 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_1 VPB VNB VGND VPWR A B Y
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211ai_1 VPB VNB VGND VPWR A1 Y C1 B1 A2
X0 a_110_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.17225 ps=1.83 w=0.65 l=0.15
X2 Y A2 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X3 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X4 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X5 a_326_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.12675 ps=1.04 w=0.65 l=0.15
X6 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.635 pd=3.27 as=0.195 ps=1.39 w=1 l=0.15
X7 Y C1 a_326_47# VNB sky130_fd_pr__nfet_01v8 ad=0.39325 pd=2.51 as=0.06825 ps=0.86 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__xnor2_1 VGND VPWR B Y A VPB VNB
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.06825 ps=0.86 w=0.65 l=0.15
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X8 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31o_2 VNB VPB VGND VPWR B1 A1 A2 A3 X
X0 VPWR A2 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1 a_277_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2 a_79_21# B1 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X3 a_277_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_361_47# A2 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_277_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12675 ps=1.04 w=0.65 l=0.15
X9 a_79_21# A1 a_361_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.10725 ps=0.98 w=0.65 l=0.15
X10 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3_2 VNB VPB VGND VPWR C A Y B
X0 VGND C a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_277_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_27_47# B a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=2.62 as=0.135 ps=1.27 w=1 l=0.15
X8 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_277_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4_2 VNB VPB VGND VPWR X D C B A
X0 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X1 VGND D a_304_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17515 pd=1.265 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.27995 ps=1.615 w=1 l=0.15
X3 a_198_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.06195 ps=0.715 w=0.42 l=0.15
X4 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X5 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X6 a_304_47# C a_198_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X7 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07455 pd=0.775 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27995 pd=1.615 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.17515 ps=1.265 w=0.65 l=0.15
X10 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.07455 ps=0.775 w=0.42 l=0.15
X11 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_2 VPWR VGND X A VPB VNB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=4.73
.ends

.subckt sky130_fd_sc_hd__a31oi_4 VNB VPB VPWR VGND Y B1 A1 A2 A3
X0 a_27_47# A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_27_47# A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.385 pd=1.77 as=0.135 ps=1.27 w=1 l=0.15
X4 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.145 ps=1.29 w=1 l=0.15
X9 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_445_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.385 ps=1.77 w=1 l=0.15
X14 a_445_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 Y A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.135 ps=1.27 w=1 l=0.15
X21 Y A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 a_445_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_445_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X28 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X31 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22o_1 VPWR VGND VPB VNB B1 A1 A2 X B2
X0 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X2 VGND A2 a_373_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X6 a_373_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X7 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X8 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux4_1 VNB VPB VGND VPWR A1 A0 S0 A3 A2 S1 X
X0 a_277_47# a_247_21# a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 VGND S0 a_247_21# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_834_97# a_247_21# a_750_97# VNB sky130_fd_pr__nfet_01v8 ad=0.10795 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VGND A3 a_668_97# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1079 ps=1.36 w=0.42 l=0.15
X4 a_1290_413# S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_834_97# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 a_750_97# S0 a_757_363# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1079 ps=1.36 w=0.42 l=0.15
X7 a_27_47# S0 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.085225 ps=0.925 w=0.42 l=0.15
X8 X a_1478_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9 VPWR A1 a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 VPWR S0 a_247_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1079 pd=1.36 as=0.1083 ps=1.36 w=0.42 l=0.15
X11 X a_1478_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X12 a_193_47# A0 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_750_97# a_1290_413# a_1478_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2688 pd=2.12 as=0.092075 ps=0.99 w=0.42 l=0.15
X14 a_1478_413# S1 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.092075 pd=0.99 as=0.1092 ps=1.36 w=0.42 l=0.15
X15 a_1290_413# S1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X16 a_277_47# a_247_21# a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.085225 pd=0.925 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 a_750_97# S0 a_668_97# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X18 a_923_363# a_247_21# a_750_97# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.090125 pd=0.995 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 a_757_363# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 VPWR A3 a_923_363# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.090125 ps=0.995 w=0.42 l=0.15
X21 a_277_47# a_1290_413# a_1478_413# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.151025 ps=1.285 w=0.42 l=0.15
X22 a_193_413# A0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X23 a_193_413# S0 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1079 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X24 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X25 a_1478_413# S1 a_750_97# VNB sky130_fd_pr__nfet_01v8 ad=0.151025 pd=1.285 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221o_1 VPWR VGND VPB VNB A1 A2 X B1 B2 C1
X0 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X2 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X5 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X6 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X7 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X9 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_4 VPWR VGND X A VPB VNB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31o_1 VPB VNB X A3 A2 A1 B1 VGND VPWR
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X1 a_209_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X2 a_303_47# A2 a_209_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X3 a_209_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X5 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X6 a_80_21# A1 a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X7 VPWR A2 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X8 a_80_21# B1 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X9 a_209_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ai_4 VNB VPB VPWR VGND B1 Y A1 A2
X0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X4 VGND A2 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X5 Y B1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6 VGND A1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X7 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 a_32_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X9 Y B1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_32_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X12 a_32_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X13 a_32_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X14 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 a_32_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.104 ps=0.97 w=0.65 l=0.15
X16 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X17 a_32_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X18 VGND A2 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X19 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X20 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X21 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X22 VGND A1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X23 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VPWR VPB VNB
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
.ends

.subckt sky130_fd_sc_hd__a211oi_1 VPWR VGND VPB VNB Y C1 B1 A1 A2
X0 a_56_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR A2 a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X3 a_139_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.2665 ps=2.12 w=0.65 l=0.15
X4 a_311_297# B1 a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X5 Y C1 a_311_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X6 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X7 Y A1 a_139_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_2 VPB VNB VPWR VGND Y A
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31a_1 X A1 A2 A3 B1 VPB VNB VGND VPWR
X0 a_103_199# B1 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X1 VPWR a_103_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
X2 a_337_297# A2 a_253_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3 a_103_199# A3 a_337_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.425 as=0.165 ps=1.33 w=1 l=0.15
X4 a_253_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X5 VPWR B1 a_103_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.2125 ps=1.425 w=1 l=0.15
X6 VGND a_103_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.234 ps=2.02 w=0.65 l=0.15
X7 a_253_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12675 ps=1.04 w=0.65 l=0.15
X8 a_253_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X9 VGND A2 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21a_1 VPB VNB VGND VPWR A1 A2 B1 X
X0 VPWR A1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X1 a_297_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X6 a_382_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a311o_1 VNB VPB VGND VPWR C1 B1 A1 A2 A3 X
X0 a_75_199# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.134875 ps=1.065 w=0.65 l=0.15
X1 a_208_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.112125 ps=0.995 w=0.65 l=0.15
X2 a_315_47# A2 a_208_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.17 as=0.125125 ps=1.035 w=0.65 l=0.15
X3 VGND B1 a_75_199# VNB sky130_fd_pr__nfet_01v8 ad=0.134875 pd=1.065 as=0.105625 ps=0.975 w=0.65 l=0.15
X4 a_75_199# A1 a_315_47# VNB sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.17 w=0.65 l=0.15
X5 a_75_199# C1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2075 ps=1.415 w=1 l=0.15
X6 a_544_297# B1 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2075 pd=1.415 as=0.1625 ps=1.325 w=1 l=0.15
X7 VPWR a_75_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.285 ps=2.57 w=1 l=0.15
X8 a_201_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1425 ps=1.285 w=1 l=0.15
X9 VPWR A2 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.165 ps=1.33 w=1 l=0.15
X10 a_201_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.305 ps=1.61 w=1 l=0.15
X11 VGND a_75_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a32o_1 VGND VPWR VPB VNB X A3 A2 A1 B1 B2
X0 a_93_21# A1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X1 a_93_21# B1 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X2 a_584_47# B1 a_93_21# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X3 VPWR a_93_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X4 VGND B2 a_584_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X5 a_256_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X6 a_250_297# B2 a_93_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 VGND a_93_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X8 a_250_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X9 VPWR A2 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X10 a_250_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X11 a_346_47# A2 a_256_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o221a_1 VPB VNB VGND VPWR B1 B2 A2 A1 X C1
X0 a_240_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_51_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VGND A1 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_51_297# B2 a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.4125 pd=1.825 as=0.105 ps=1.21 w=1 l=0.15
X4 a_149_47# C1 a_51_297# VNB sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.2015 ps=1.92 w=0.65 l=0.15
X5 a_240_47# B1 a_149_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.099125 ps=0.955 w=0.65 l=0.15
X6 VPWR A1 a_512_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X7 X a_51_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.165 ps=1.33 w=1 l=0.15
X8 a_149_47# B2 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_245_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X10 VPWR C1 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.34 ps=2.68 w=1 l=0.15
X11 a_512_297# A2 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.4125 ps=1.825 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_8 X A VPB VNB VGND VPWR
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X11 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X18 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4b_1 VPWR VGND VPB VNB B C A X D_N
X0 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X1 a_109_53# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_215_297# a_109_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.101875 ps=0.99 w=0.65 l=0.15
X4 a_392_297# C a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.04515 pd=0.635 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 a_465_297# B a_392_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06405 pd=0.725 as=0.04515 ps=0.635 w=0.42 l=0.15
X6 a_215_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VPWR A a_465_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06405 ps=0.725 w=0.42 l=0.15
X8 a_297_297# a_109_53# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_109_53# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 VGND C a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06405 ps=0.725 w=0.42 l=0.15
X11 VGND A a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ba_1 VNB VPB VGND VPWR B1_N A1 A2 X
X0 a_222_93# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X1 VPWR A1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X2 VGND a_79_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_222_93# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.18575 ps=1.415 w=0.42 l=0.15
X4 VGND A2 a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X5 a_448_47# a_222_93# a_79_199# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_79_199# a_222_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X7 a_544_297# A2 a_79_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X8 a_448_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR a_79_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18575 pd=1.415 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 VNB VPB VGND VPWR A X
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21bo_1 VNB VPB VGND VPWR X A2 A1 B1_N
X0 a_298_297# a_27_413# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1 a_215_297# a_27_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1359 ps=1.1 w=0.65 l=0.15
X2 a_298_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.258375 ps=1.445 w=0.65 l=0.15
X4 VPWR B1_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6 a_382_47# A1 a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND B1_N a_27_413# VNB sky130_fd_pr__nfet_01v8 ad=0.1359 pd=1.1 as=0.1113 ps=1.37 w=0.42 l=0.15
X8 VPWR A1 a_298_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND A2 a_382_47# VNB sky130_fd_pr__nfet_01v8 ad=0.258375 pd=1.445 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2b_1 X A_N B VGND VPWR VPB VNB
X0 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X2 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o41a_1 VPB VNB VGND VPWR X B1 A4 A3 A2 A1
X0 VGND A4 a_321_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_321_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.1235 ps=1.03 w=0.65 l=0.15
X2 a_103_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=1.52 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR a_103_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.425 ps=2.85 w=1 l=0.15
X4 VGND a_103_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.247 ps=2.06 w=0.65 l=0.15
X5 VGND A2 a_321_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X6 a_321_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.12675 ps=1.04 w=0.65 l=0.15
X7 a_511_297# A3 a_393_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.22 ps=1.44 w=1 l=0.15
X8 a_619_297# A2 a_511_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X9 a_321_47# B1 a_103_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 a_393_297# A4 a_103_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.26 ps=1.52 w=1 l=0.15
X11 VPWR A1 a_619_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.195 ps=1.39 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4_1 X C A B D VGND VPWR VPB VNB
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_4 VPB VNB VGND VPWR Y B A
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X11 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_1 VPWR VGND VPB VNB B C A X
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.101875 ps=0.99 w=0.65 l=0.15
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3b_1 A_N B X C VGND VPWR VPB VNB
X0 a_109_93# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 X a_209_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X2 a_109_93# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 a_296_53# a_109_93# a_209_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X4 VPWR C a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X5 a_368_53# B a_296_53# VNB sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_209_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
X7 a_209_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VPWR a_109_93# a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X9 VGND C a_368_53# VNB sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2_2 VPWR VGND A X B VPB VNB
X0 X a_61_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.16655 ps=1.39 w=1 l=0.15
X1 VPWR a_61_75# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X2 VPWR B a_61_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VGND B a_147_75# VNB sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 X a_61_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.1118 ps=1.04 w=0.65 l=0.15
X5 VGND a_61_75# X VNB sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X6 a_61_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X7 a_147_75# A a_61_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 VGND VPWR A X VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_2 VPWR VGND VPB VNB X A B
X0 a_121_297# B a_39_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 X a_39_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10675 ps=1.005 w=0.65 l=0.15
X2 VPWR a_39_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_39_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15575 ps=1.355 w=1 l=0.15
X4 VGND a_39_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR A a_121_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15575 pd=1.355 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VGND A a_39_297# VNB sky130_fd_pr__nfet_01v8 ad=0.10675 pd=1.005 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_39_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux2_4 VNB VPB VPWR VGND X S A1 A0
X0 a_204_297# A1 a_396_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.16 ps=1.32 w=1 l=0.15
X1 VPWR a_396_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 X a_396_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR S a_314_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 a_204_297# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1625 ps=1.325 w=1 l=0.15
X5 a_396_47# A0 a_314_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.26 ps=2.52 w=1 l=0.15
X6 a_206_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.108875 ps=0.985 w=0.65 l=0.15
X7 X a_396_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 X a_396_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR a_396_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 a_490_47# A1 a_396_47# VNB sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.104 ps=0.97 w=0.65 l=0.15
X11 VGND S a_490_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.274625 ps=1.495 w=0.65 l=0.15
X12 VGND a_396_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_396_47# A0 a_206_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.26 ps=1.45 w=0.65 l=0.15
X14 VGND a_396_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VPWR S a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X16 X a_396_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND S a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.108875 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_1 VGND VPWR X A VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3_1 VPB VNB VGND VPWR C B A Y
X0 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_109_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22o_4 VNB VPB VGND VPWR X B2 A1 A2 B1
X0 a_484_297# B2 a_96_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND B2 a_566_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 X a_96_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VPWR a_96_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_96_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_96_21# B1 a_484_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR a_96_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 X a_96_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X8 VGND a_96_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_484_297# B1 a_96_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_484_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND A2 a_918_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_96_21# B2 a_484_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 a_96_21# B1 a_566_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_484_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VPWR A1 a_484_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_96_21# A1 a_918_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VPWR A2 a_484_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X18 a_566_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25675 ps=1.44 w=0.65 l=0.15
X19 a_918_47# A1 a_96_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_566_47# B1 a_96_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 a_918_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X22 X a_96_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X23 VGND a_96_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 VPWR VGND VPB VNB X A
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22a_1 VPB VNB VGND VPWR B2 A2 A1 B1 X
X0 a_78_199# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2 a_493_297# A2 a_78_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X3 VPWR a_78_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3725 pd=1.745 as=0.28 ps=2.56 w=1 l=0.15
X4 VGND A2 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X5 a_78_199# B2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.1175 ps=1.235 w=1 l=0.15
X6 a_215_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_215_47# B2 a_78_199# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_292_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1175 pd=1.235 as=0.3725 ps=1.745 w=1 l=0.15
X9 VGND a_78_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_1 VPWR VGND VPB VNB B D C A X
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211ai_2 VNB VPB VGND VPWR Y B1 A2 A1 C1
X0 a_286_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2 a_286_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X3 Y A2 a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4 VGND A1 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X5 Y C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X6 VGND A2 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X7 a_487_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 a_27_47# B1 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10 VPWR A1 a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_27_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X12 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X13 a_487_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X14 a_286_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X15 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4bb_2 VNB VPB VGND VPWR A_N X C D B_N
X0 a_174_21# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1 a_174_21# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.33075 ps=1.705 w=0.42 l=0.15
X2 a_476_47# a_27_47# a_174_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.33075 pd=1.705 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14075 ps=1.325 w=1 l=0.15
X5 a_548_47# a_505_280# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X8 VPWR D a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 VGND D a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 VPWR a_505_280# a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X11 a_505_280# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0924 ps=0.86 w=0.42 l=0.15
X12 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_505_280# B_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0924 ps=0.86 w=0.42 l=0.15
X14 a_639_47# C a_548_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06405 ps=0.725 w=0.42 l=0.15
X15 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_2 VPB VNB VGND VPWR Y A B
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3_2 B X A C VPWR VGND VPB VNB
X0 VPWR a_29_311# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_29_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15075 ps=1.345 w=1 l=0.15
X2 VPWR A a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND a_29_311# X VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_184_53# B a_112_53# VNB sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X5 VPWR C a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15075 pd=1.345 as=0.074375 ps=0.815 w=0.42 l=0.15
X6 X a_29_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1304 ps=1.105 w=0.65 l=0.15
X7 a_112_53# A a_29_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_29_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 VGND C a_184_53# VNB sky130_fd_pr__nfet_01v8 ad=0.1304 pd=1.105 as=0.05355 ps=0.675 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3_1 VPB VNB VGND VPWR A B Y C
X0 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X2 a_193_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X4 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 a_109_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_4 VNB VPB VGND VPWR B A X
X0 a_121_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X1 VPWR a_35_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2 X a_35_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_35_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X4 X a_35_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR a_35_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 X a_35_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X7 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR A a_121_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X9 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfxtp_4 VGND VPWR VNB VPB Q D CLK
X0 Q a_1062_300# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1425 ps=1.285 w=1 l=0.15
X1 a_1020_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0657 ps=0.725 w=0.36 l=0.15
X2 a_572_47# a_193_47# a_475_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0687 pd=0.76 as=0.0594 ps=0.69 w=0.36 l=0.15
X3 VPWR a_1062_300# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1218 pd=1.42 as=0.09135 ps=0.855 w=0.42 l=0.15
X4 a_634_183# a_475_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.1493 ps=1.22 w=0.64 l=0.15
X5 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 a_475_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X8 VGND a_1062_300# a_1020_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1197 pd=1.41 as=0.066 ps=0.745 w=0.42 l=0.15
X9 VPWR a_634_183# a_568_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 Q a_1062_300# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.092625 ps=0.935 w=0.65 l=0.15
X11 a_568_413# a_27_47# a_475_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.06615 ps=0.735 w=0.42 l=0.15
X12 a_634_183# a_475_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X13 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.09135 pd=0.855 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_891_413# a_27_47# a_634_183# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X16 Q a_1062_300# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.105625 ps=0.975 w=0.65 l=0.15
X17 VGND a_891_413# a_1062_300# VNB sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X18 VPWR a_1062_300# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.135 ps=1.27 w=1 l=0.15
X19 VGND a_1062_300# Q VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 Q a_1062_300# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X22 VGND a_1062_300# Q VNB sky130_fd_pr__nfet_01v8 ad=0.092625 pd=0.935 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X24 VPWR a_891_413# a_1062_300# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.28 ps=2.56 w=1 l=0.15
X25 a_891_413# a_193_47# a_634_183# VNB sky130_fd_pr__nfet_01v8 ad=0.0657 pd=0.725 as=0.0989 ps=0.995 w=0.36 l=0.15
X26 a_475_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0672 ps=0.74 w=0.42 l=0.15
X27 VGND a_634_183# a_572_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1493 pd=1.22 as=0.0687 ps=0.76 w=0.42 l=0.15
X28 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X29 VPWR a_1062_300# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2b_2 VPWR VGND VNB VPB A B_N X
X0 VPWR A a_300_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_218_297# a_27_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.15645 ps=1.165 w=0.42 l=0.15
X2 VGND B_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0.15645 pd=1.165 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 a_300_297# a_27_53# a_218_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 X a_218_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.101875 ps=0.99 w=0.65 l=0.15
X5 VPWR a_218_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=2.62 as=0.135 ps=1.27 w=1 l=0.15
X6 X a_218_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14825 ps=1.34 w=1 l=0.15
X7 VGND a_218_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_27_53# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 VGND A a_218_297# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21boi_1 VPWR VGND VPB VNB B1_N Y A1 A2
X0 a_300_297# a_27_413# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR B1_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.15
X3 Y a_27_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.101875 ps=0.99 w=0.65 l=0.15
X4 VPWR A1 a_300_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 a_384_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.143 ps=1.09 w=0.65 l=0.15
X6 VGND B1_N a_27_413# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.1113 ps=1.37 w=0.42 l=0.15
X7 a_300_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ai_2 VGND VPWR B1 A1 Y A2 VPB VNB
X0 VGND A2 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X1 Y B1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 VPWR A1 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.175 ps=1.35 w=1 l=0.15
X4 a_29_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5 Y A2 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND A1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X7 a_112_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X8 a_112_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.14 ps=1.28 w=1 l=0.15
X9 a_29_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X11 a_29_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.12675 ps=1.04 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3_4 VPB VNB VGND VPWR B A Y C
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_449_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_27_297# B a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 Y C a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_449_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y C a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X10 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_449_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X15 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_27_297# B a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 a_449_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4bb_1 VNB VPB VGND VPWR A_N B_N C D X
X0 VPWR D a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.46 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_223_47# B_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1386 pd=1.5 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 a_515_93# a_223_47# a_429_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 a_223_47# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1344 pd=1.48 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X5 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X6 X a_343_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.172 ps=1.46 w=1 l=0.15
X7 a_429_93# a_27_47# a_343_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1176 ps=1.4 w=0.42 l=0.15
X8 VGND D a_615_93# VNB sky130_fd_pr__nfet_01v8 ad=0.1265 pd=1.11 as=0.0777 ps=0.79 w=0.42 l=0.15
X9 a_343_93# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X10 a_343_93# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X11 a_615_93# C a_515_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X12 X a_343_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1654 pd=1.82 as=0.1265 ps=1.11 w=0.65 l=0.15
X13 VPWR a_223_47# a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3b_2 VPWR VGND VPB VNB C_N X A B
X0 a_388_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.14825 ps=1.34 w=0.42 l=0.15
X1 VPWR C_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X4 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X7 a_176_21# a_27_47# a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 a_472_297# B a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.101875 ps=0.99 w=0.42 l=0.15
X10 a_176_21# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 VGND C_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2bb2a_1 VNB VPB VPWR VGND X A1_N A2_N B2 B1
X0 a_206_369# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.14575 ps=1.335 w=0.42 l=0.15
X1 a_206_369# A2_N a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06615 ps=0.735 w=0.42 l=0.15
X2 VGND B2 a_489_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_585_369# B2 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0672 ps=0.74 w=0.42 l=0.15
X4 a_489_47# a_206_369# a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_489_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VPWR A2_N a_206_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.20925 pd=1.345 as=0.129 ps=1.18 w=0.42 l=0.15
X7 a_76_199# a_206_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.20925 ps=1.345 w=0.42 l=0.15
X8 a_205_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06615 pd=0.735 as=0.098625 ps=0.98 w=0.42 l=0.15
X9 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X10 VPWR B1 a_585_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.098625 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_4 VNB VPB VPWR VGND D C B A X
X0 VPWR A a_304_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X1 a_304_297# B a_220_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND C a_32_297# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X3 a_220_297# C a_114_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X4 a_32_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_32_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR a_32_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X7 X a_32_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND A a_32_297# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR a_32_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 X a_32_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X11 X a_32_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 X a_32_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X13 a_114_297# D a_32_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.26 ps=2.52 w=1 l=0.15
X14 VGND a_32_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VGND a_32_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2111a_1 VNB VPB VPWR VGND X D1 C1 B1 A2 A1
X0 a_676_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.2125 ps=1.425 w=1 l=0.15
X1 a_512_47# B1 a_409_47# VNB sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.118625 ps=1.015 w=0.65 l=0.15
X2 a_306_47# D1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.19825 ps=1.91 w=0.65 l=0.15
X3 VGND A2 a_512_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.19825 ps=1.26 w=0.65 l=0.15
X4 VPWR C1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.2175 ps=1.435 w=1 l=0.15
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.425 as=0.305 ps=1.61 w=1 l=0.15
X6 VPWR A1 a_676_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X7 a_512_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_409_47# C1 a_306_47# VNB sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.118625 ps=1.015 w=0.65 l=0.15
X9 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3825 pd=1.765 as=0.26 ps=2.52 w=1 l=0.15
X10 a_79_21# D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2175 pd=1.435 as=0.3825 ps=1.765 w=1 l=0.15
X11 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21bai_1 VPB VNB VPWR VGND A1 B1_N Y A2
X0 a_388_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1275 pd=1.255 as=0.1525 ps=1.305 w=1 l=0.15
X1 a_105_352# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_297_47# a_105_352# Y VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR A1 a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1275 ps=1.255 w=1 l=0.15
X5 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X6 VPWR B1_N a_105_352# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17825 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 Y a_105_352# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.17825 ps=1.4 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2b_2 VPB VNB VGND VPWR Y A B_N
X0 Y a_251_21# a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y a_251_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17875 ps=1.85 w=0.65 l=0.15
X5 VGND a_251_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7 VPWR B_N a_251_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 VGND B_N a_251_21# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_27_297# a_251_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_2 VGND VPWR VPB VNB B C A X
X0 VPWR a_30_53# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.315 pd=2.63 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND a_30_53# X VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 X a_30_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14825 ps=1.34 w=1 l=0.15
X3 a_112_297# C a_30_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 X a_30_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.101875 ps=0.99 w=0.65 l=0.15
X5 VGND A a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 a_30_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VGND C a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_184_297# B a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X9 VPWR A a_184_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a41o_1 VGND VPWR A3 A4 A2 X B1 A1 VPB VNB
X0 a_465_47# A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VGND A4 a_561_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 VPWR A3 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3 a_297_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4 a_297_297# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X5 VPWR A1 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_381_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.183625 ps=1.215 w=0.65 l=0.15
X7 a_297_297# B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X9 a_79_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.183625 pd=1.215 as=0.160875 ps=1.145 w=0.65 l=0.15
X10 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.160875 pd=1.145 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_561_47# A3 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__xor2_2 VPWR VGND X B A VPB VNB
X0 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_470_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_470_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR A a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_470_47# B X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.105625 ps=0.975 w=0.65 l=0.15
X6 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17875 ps=1.85 w=0.65 l=0.15
X8 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.275 ps=2.55 w=1 l=0.15
X10 a_470_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1625 ps=1.325 w=1 l=0.15
X11 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12 VPWR B a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X13 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VGND A a_470_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X16 X a_112_47# a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 a_470_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X18 X B a_470_47# VNB sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4b_4 VNB VPB VGND VPWR X D_N C B A
X0 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND a_215_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VPWR a_215_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_109_93# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 a_215_297# a_109_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.16535 ps=1.82 w=0.65 l=0.15
X5 VGND C a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X6 VGND A a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X8 a_215_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_109_93# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 VPWR A a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND a_215_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_487_297# B a_403_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_403_297# C a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X14 VPWR a_215_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X16 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_297_297# a_109_93# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4bb_4 VNB VPB VGND VPWR B A X C_N D_N
X0 VPWR a_315_380# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_315_380# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X2 a_315_380# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND C_N a_27_410# VNB sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VPWR C_N a_27_410# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1226 pd=1.32 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VPWR A a_583_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND a_27_410# a_315_380# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X7 a_583_297# B a_499_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND A a_315_380# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_397_297# a_205_93# a_315_380# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.257925 ps=2.52 w=1 l=0.15
X10 X a_315_380# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X11 X a_315_380# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_499_297# a_27_410# a_397_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.18 ps=1.36 w=1 l=0.15
X13 VPWR a_315_380# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14 a_205_93# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06195 ps=0.715 w=0.42 l=0.15
X15 a_205_93# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11295 pd=1.4 as=0.1226 ps=1.32 w=0.42 l=0.15
X16 VGND a_315_380# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VGND a_315_380# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_315_380# a_205_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.169 ps=1.82 w=0.65 l=0.15
X19 X a_315_380# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_2 VNB VPB VGND VPWR A2 A1 Y B1
X0 VGND A2 a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X1 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=2.1 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y A1 a_114_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X3 a_114_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.18525 ps=1.87 w=0.65 l=0.15
X4 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X8 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X10 a_285_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.091 ps=0.93 w=0.65 l=0.15
X11 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22ai_1 VPB VNB VGND VPWR A1 A2 B1 B2 Y
X0 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X1 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.092625 ps=0.935 w=0.65 l=0.15
X2 VPWR A1 a_307_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.105 ps=1.21 w=1 l=0.15
X3 a_307_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.2325 ps=1.465 w=1 l=0.15
X4 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2325 pd=1.465 as=0.1125 ps=1.225 w=1 l=0.15
X6 a_109_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1125 pd=1.225 as=0.26 ps=2.52 w=1 l=0.15
X7 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.092625 pd=0.935 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4_4 VNB VPB VGND VPWR X D C B A
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_188_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.108875 pd=0.985 as=0.079625 ps=0.895 w=0.65 l=0.15
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND D a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.141375 ps=1.085 w=0.65 l=0.15
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.215 ps=1.43 w=1 l=0.15
X6 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.135 ps=1.27 w=1 l=0.15
X9 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.105625 ps=0.975 w=0.65 l=0.15
X10 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.215 pd=1.43 as=0.155 ps=1.31 w=1 l=0.15
X12 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X14 a_285_47# C a_188_47# VNB sky130_fd_pr__nfet_01v8 ad=0.141375 pd=1.085 as=0.108875 ps=0.985 w=0.65 l=0.15
X15 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.079625 pd=0.895 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2bb2o_1 VNB VPB VGND VPWR B1 A1_N A2_N X B2
X0 a_226_47# A2_N a_226_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_489_413# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_226_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.16675 ps=1.435 w=0.42 l=0.15
X3 VPWR B2 a_489_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_489_413# a_226_47# a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_76_199# a_226_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1386 ps=1.08 w=0.42 l=0.15
X6 VGND B1 a_556_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_556_47# B2 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND A2_N a_226_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1386 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_226_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1201 ps=1.085 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16675 pd=1.435 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.1201 pd=1.085 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2111oi_1 VNB VPWR VGND VPB D1 C1 B1 A1 Y A2
X0 a_316_297# C1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.1725 ps=1.345 w=1 l=0.15
X1 Y D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.481 ps=2.78 w=0.65 l=0.15
X2 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.12025 pd=1.02 as=0.125125 ps=1.035 w=0.65 l=0.15
X3 a_420_297# B1 a_316_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=1.58 as=0.185 ps=1.37 w=1 l=0.15
X4 VPWR A1 a_420_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.29 ps=1.58 w=1 l=0.15
X5 VGND A2 a_568_47# VNB sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.89 as=0.0845 ps=0.91 w=0.65 l=0.15
X6 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.24 as=0.12025 ps=1.02 w=0.65 l=0.15
X7 a_420_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.1375 ps=1.275 w=1 l=0.15
X8 a_217_297# D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.755 ps=3.51 w=1 l=0.15
X9 a_568_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0845 pd=0.91 as=0.19175 ps=1.24 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o221a_2 VPB VNB VGND VPWR B1 B2 A2 A1 X C1
X0 VPWR a_38_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR A1 a_497_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X2 X a_38_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X3 a_141_47# B2 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_497_297# A2 a_38_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.3875 ps=1.775 w=1 l=0.15
X5 VGND A1 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR C1 a_38_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.325 ps=2.65 w=1 l=0.15
X7 a_237_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1125 pd=1.225 as=0.165 ps=1.33 w=1 l=0.15
X8 a_38_47# B2 a_237_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3875 pd=1.775 as=0.1125 ps=1.225 w=1 l=0.15
X9 a_225_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 X a_38_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_141_47# C1 a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.23725 ps=2.03 w=0.65 l=0.15
X12 VGND a_38_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_225_47# B1 a_141_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_4 VPB VNB VPWR VGND B C A X
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.26 ps=1.45 w=0.65 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.4 ps=1.8 w=1 l=0.15
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.20475 pd=1.93 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.4 pd=1.8 as=0.135 ps=1.27 w=1 l=0.15
X5 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_109_297# C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 VGND C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2111o_1 VPB VGND VPWR VNB B1 X D1 A1 A2 C1
X0 VGND A2 a_660_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X1 VGND C1 a_85_193# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X2 a_414_297# C1 a_334_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X3 VGND a_85_193# X VNB sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X4 a_334_297# D1 a_85_193# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X5 a_516_297# B1 a_414_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X6 a_516_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X7 a_660_47# A1 a_85_193# VNB sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X8 a_85_193# D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X9 VPWR A1 a_516_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X10 a_85_193# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X11 VPWR a_85_193# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2111o_2 VNB VPB VGND VPWR A2 A1 B1 C1 X D1
X0 VPWR a_86_235# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1 VGND C1 a_86_235# VNB sky130_fd_pr__nfet_01v8 ad=0.121875 pd=1.025 as=0.091 ps=0.93 w=0.65 l=0.15
X2 X a_86_235# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 a_86_235# D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.290875 ps=1.545 w=0.65 l=0.15
X4 X a_86_235# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X5 a_715_47# A1 a_86_235# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.108875 ps=0.985 w=0.65 l=0.15
X6 VGND A2 a_715_47# VNB sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.12675 ps=1.04 w=0.65 l=0.15
X7 a_499_297# C1 a_427_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X8 VGND a_86_235# X VNB sky130_fd_pr__nfet_01v8 ad=0.290875 pd=1.545 as=0.091 ps=0.93 w=0.65 l=0.15
X9 a_86_235# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.108875 pd=0.985 as=0.121875 ps=1.025 w=0.65 l=0.15
X10 a_607_297# B1 a_499_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X11 a_427_297# D1 a_86_235# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.41 ps=2.82 w=1 l=0.15
X12 VPWR A1 a_607_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X13 a_607_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.195 ps=1.39 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21bai_2 VNB VPB VGND VPWR B1_N Y A2 A1
X0 a_397_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR B1_N a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 Y A2 a_397_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3 VGND A2 a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VGND A1 a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_28_297# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 Y a_28_297# a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 VPWR a_28_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8 a_397_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X9 a_229_47# a_28_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y a_28_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X11 a_229_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_229_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VPWR A1 a_397_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4b_2 VPWR VGND VPB VNB C D_N X A B
X0 a_176_21# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 VGND D_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X4 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16835 pd=1.495 as=0.135 ps=1.27 w=1 l=0.15
X5 a_555_297# C a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 a_176_21# a_27_53# a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1693 ps=1.5 w=1 l=0.15
X8 a_387_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.16835 ps=1.495 w=0.42 l=0.15
X9 a_483_297# B a_387_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 VGND a_27_53# a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 VPWR D_N a_27_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1693 pd=1.5 as=0.1092 ps=1.36 w=0.42 l=0.15
X13 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.10025 ps=0.985 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3b_1 VPB VNB VGND VPWR Y B C A_N
X0 Y a_53_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1925 ps=1.385 w=1 l=0.15
X1 a_232_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR A_N a_53_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VGND A_N a_53_93# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_316_47# B a_232_47# VNB sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y a_53_93# a_316_47# VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.125125 ps=1.035 w=0.65 l=0.15
X7 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__xnor2_4 VNB VPB VGND VPWR Y B A
X0 VGND A a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 Y a_38_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_38_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_820_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR a_38_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X5 VGND A a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VGND B a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND B a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y B a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_38_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 a_38_297# B a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VGND A a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_902_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_820_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 a_902_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VPWR A a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 Y a_38_297# a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X17 Y a_38_297# a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_38_47# B a_38_297# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_38_47# B a_38_297# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_38_297# B a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X21 a_38_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 VPWR B a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X23 a_38_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 a_902_47# a_38_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 a_902_47# a_38_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 Y B a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_38_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 a_820_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 VPWR A a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 VGND A a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 VPWR A a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 a_902_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X33 a_820_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 Y a_38_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X35 a_902_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X36 a_38_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 VPWR A a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X38 VPWR a_38_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X39 VPWR B a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o311a_1 X A1 A2 A3 B1 C1 VPB VNB VGND VPWR
X0 a_585_47# B1 a_266_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.118625 ps=1.015 w=0.65 l=0.15
X1 VGND A2 a_266_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.07 as=0.117 ps=1.01 w=0.65 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3125 pd=1.625 as=0.26 ps=2.52 w=1 l=0.15
X3 a_81_21# C1 a_585_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.203125 pd=1.275 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_266_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.3125 ps=1.625 w=1 l=0.15
X6 a_368_297# A2 a_266_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.18 ps=1.36 w=1 l=0.15
X7 a_266_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.1365 ps=1.07 w=0.65 l=0.15
X8 a_266_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.203125 ps=1.275 w=0.65 l=0.15
X9 a_81_21# A3 a_368_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.21 ps=1.42 w=1 l=0.15
X10 a_81_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X11 VPWR B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.1375 ps=1.275 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a32o_2 VNB VPB VGND VPWR X A3 A2 B2 B1 A1
X0 VPWR A3 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.215 ps=1.43 w=1 l=0.15
X2 a_352_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.209625 ps=1.295 w=0.65 l=0.15
X3 a_549_47# A1 a_21_199# VNB sky130_fd_pr__nfet_01v8 ad=0.13975 pd=1.08 as=0.10725 ps=0.98 w=0.65 l=0.15
X4 X a_21_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND a_21_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.209625 pd=1.295 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_665_47# A2 a_549_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13975 ps=1.08 w=0.65 l=0.15
X7 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.215 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X8 a_299_297# B1 a_21_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_21_199# B2 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 VGND A3 a_665_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VPWR a_21_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 X a_21_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_21_199# B1 a_352_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.115375 ps=1.005 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31a_4 VGND VPWR VPB VNB X A2 A1 A3 B1
X0 VPWR A1 a_926_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND A1 a_496_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_926_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A3 a_496_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X4 VGND a_102_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND A2 a_496_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_926_297# A2 a_672_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_102_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.135 ps=1.27 w=1 l=0.15
X8 a_496_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 X a_102_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.0975 ps=0.95 w=0.65 l=0.15
X10 a_102_21# B1 a_496_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X11 VPWR a_102_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 X a_102_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 X a_102_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15 ps=1.3 w=1 l=0.15
X14 VPWR a_102_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.135 ps=1.27 w=1 l=0.15
X15 a_672_297# A3 a_102_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_496_47# B1 a_102_21# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_102_21# A3 a_672_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X18 VGND a_102_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 X a_102_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X20 a_496_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 VPWR B1 a_102_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.145 ps=1.29 w=1 l=0.15
X22 a_496_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 a_672_297# A2 a_926_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__xnor2_2 VGND VPWR Y A B VPB VNB
X0 a_27_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_560_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2 VGND B a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.099125 ps=0.955 w=0.65 l=0.15
X3 Y B a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y a_27_297# a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_474_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X7 VGND A a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_27_47# B a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_27_297# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17875 ps=1.85 w=0.65 l=0.15
X10 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VPWR B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.275 ps=2.55 w=1 l=0.15
X12 a_474_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_560_47# a_27_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14 VPWR A a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X15 Y a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X16 VPWR a_27_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X17 a_560_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211o_2 VNB VPB VGND VPWR X A2 A1 B1 C1
X0 a_79_21# A1 a_348_47# VNB sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.13325 ps=1.06 w=0.65 l=0.15
X1 a_79_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.199875 pd=1.265 as=0.091 ps=0.93 w=0.65 l=0.15
X3 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 a_79_21# C1 a_585_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5 VPWR A2 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X6 a_299_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.195 ps=1.39 w=1 l=0.15
X7 a_585_297# B1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X8 a_348_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.13325 pd=1.06 as=0.199875 ps=1.265 w=0.65 l=0.15
X9 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.115375 ps=1.005 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2b_1 VGND VPWR VNB VPB A X B_N
X0 a_219_297# a_27_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1575 ps=1.17 w=0.42 l=0.15
X1 VGND B_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.17 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VPWR A a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 X a_219_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X4 a_301_297# a_27_53# a_219_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 X a_219_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X6 a_27_53# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 VGND A a_219_297# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux4_2 VNB VPB VGND VPWR S0 A2 A3 S1 A1 A0 X
X0 a_600_345# S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1 a_788_316# S1 a_288_47# VNB sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VPWR A3 a_372_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1645 ps=1.33 w=0.64 l=0.15
X3 a_872_316# a_600_345# a_788_316# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X4 VPWR S0 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5 a_1279_413# S0 a_872_316# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.10535 pd=0.995 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND a_788_316# X VNB sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_1060_369# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.13775 pd=1.165 as=0.1664 ps=1.8 w=0.64 l=0.15
X8 a_872_316# a_27_47# a_1060_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.13775 ps=1.165 w=0.42 l=0.15
X9 a_1281_47# a_27_47# a_872_316# VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.072 ps=0.76 w=0.36 l=0.15
X10 a_193_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 a_1064_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0786 pd=0.805 as=0.1092 ps=1.36 w=0.42 l=0.15
X12 a_872_316# S1 a_788_316# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1404 pd=1.6 as=0.0729 ps=0.81 w=0.54 l=0.15
X13 a_872_316# S0 a_1064_47# VNB sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.0786 ps=0.805 w=0.36 l=0.15
X14 X a_788_316# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10675 ps=1.005 w=0.65 l=0.15
X15 a_788_316# a_600_345# a_288_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0729 pd=0.81 as=0.1404 ps=1.6 w=0.54 l=0.15
X16 a_372_413# a_27_47# a_288_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1645 pd=1.33 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 VGND A3 a_397_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.06705 ps=0.75 w=0.42 l=0.15
X18 a_600_345# S1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0.0819 ps=0.81 w=0.42 l=0.15
X19 a_193_369# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.09575 pd=0.965 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 VPWR a_788_316# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.135 ps=1.27 w=1 l=0.15
X21 a_288_47# S0 a_193_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.09575 ps=0.965 w=0.42 l=0.15
X22 a_397_47# S0 a_288_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06705 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X23 VGND A0 a_1281_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10675 pd=1.005 as=0.066 ps=0.745 w=0.42 l=0.15
X24 a_288_47# a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X25 X a_788_316# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.154 ps=1.335 w=1 l=0.15
X26 VGND S0 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X27 VPWR A0 a_1279_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.10535 ps=0.995 w=0.64 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22a_2 VNB VPB VGND VPWR A1 A2 B2 B1 X
X0 a_301_47# B2 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VGND A2 a_301_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X2 a_383_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.39 ps=1.78 w=1 l=0.15
X3 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.39 pd=1.78 as=0.135 ps=1.27 w=1 l=0.15
X4 a_301_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 X a_81_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 X a_81_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X8 VPWR A1 a_579_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X9 a_81_21# B1 a_301_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 a_579_297# A2 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X11 a_81_21# B2 a_383_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.105 ps=1.21 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21o_2 VNB VPB VGND VPWR A2 A1 B1 X
X0 VPWR a_80_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1 X a_80_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 VGND a_80_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.1105 pd=0.99 as=0.091 ps=0.93 w=0.65 l=0.15
X3 a_386_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X4 X a_80_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X5 a_80_199# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1625 pd=1.15 as=0.1105 ps=0.99 w=0.65 l=0.15
X6 a_386_297# B1 a_80_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_458_47# A1 a_80_199# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.1625 ps=1.15 w=0.65 l=0.15
X8 VPWR A1 a_386_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.14 ps=1.28 w=1 l=0.15
X9 VGND A2 a_458_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.1235 ps=1.03 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21boi_2 VNB VPB VPWR VGND B1_N A2 Y A1
X0 Y a_61_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.183125 ps=1.24 w=0.65 l=0.15
X1 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_217_297# a_61_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_479_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X4 a_217_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X5 Y a_61_47# a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VPWR A1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_61_47# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.15
X8 VGND A2 a_637_47# VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND a_61_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y A1 a_479_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.06825 ps=0.86 w=0.65 l=0.15
X11 VGND B1_N a_61_47# VNB sky130_fd_pr__nfet_01v8 ad=0.183125 pd=1.24 as=0.126 ps=1.44 w=0.42 l=0.15
X12 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X13 a_637_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21bai_4 VNB VPB VGND VPWR A2 A1 B1_N Y
X0 Y a_33_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_225_47# a_33_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VPWR a_33_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_33_297# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.182 ps=1.86 w=0.65 l=0.15
X4 Y a_33_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A2 a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 Y a_33_297# a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 Y a_33_297# a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VGND A2 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VGND A2 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 a_561_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X11 a_225_47# a_33_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VPWR A1 a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_225_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_225_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_225_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_225_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VPWR A1 a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 a_561_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR B1_N a_33_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X20 a_561_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 VGND A1 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 Y A2 a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VGND A1 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 a_561_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 VPWR a_33_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor4b_2 VNB VPB VGND VPWR A B C Y D_N
X0 VPWR D_N a_694_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 a_27_297# B a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_474_297# a_694_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_277_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 Y a_694_21# a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VGND D_N a_694_21# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_474_297# C a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 Y a_694_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_277_297# C a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND a_694_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21o_4 VNB VPB VGND VPWR X B1 A1 A2
X0 VGND B1 a_84_21# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_741_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X2 a_84_21# A1 a_741_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.07475 ps=0.88 w=0.65 l=0.15
X3 VGND A2 a_901_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR a_84_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR A2 a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_483_297# B1 a_84_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 X a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X8 a_84_21# B1 a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VGND a_84_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.264875 pd=1.465 as=0.091 ps=0.93 w=0.65 l=0.15
X10 VPWR a_84_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_483_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=2.79 as=0.135 ps=1.27 w=1 l=0.15
X12 VPWR A1 a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 VGND a_84_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X14 X a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.285 ps=2.57 w=1 l=0.15
X15 a_84_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.264875 ps=1.465 w=0.65 l=0.15
X16 a_483_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 X a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X18 a_901_47# A1 a_84_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 X a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31o_4 VNB VPB VGND VPWR X B1 A2 A1 A3
X0 VPWR a_277_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_277_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 X a_277_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X5 a_277_47# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X6 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND a_277_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND a_277_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_193_47# A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_361_47# A1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 X a_277_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VGND A3 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X15 X a_277_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25675 ps=1.44 w=0.65 l=0.15
X16 a_277_47# A1 a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_445_47# A2 a_361_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VGND B1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_27_297# B1 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X21 VPWR a_277_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.5 pd=3 as=0.135 ps=1.27 w=1 l=0.15
X22 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X23 a_277_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4b_2 VPWR VGND VNB VPB A_N B C D X
X0 VPWR a_193_413# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X1 a_297_47# a_27_413# a_193_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_369_47# B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 X a_193_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.103975 ps=1 w=0.65 l=0.15
X4 VPWR D a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14325 pd=1.33 as=0.06615 ps=0.735 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VGND D a_469_47# VNB sky130_fd_pr__nfet_01v8 ad=0.103975 pd=1 as=0.06195 ps=0.715 w=0.42 l=0.15
X7 VGND a_193_413# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.099125 ps=0.955 w=0.65 l=0.15
X8 VPWR B a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X9 a_193_413# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.1281 ps=1.03 w=0.42 l=0.15
X10 X a_193_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.14325 ps=1.33 w=1 l=0.15
X11 a_193_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 a_469_47# C a_369_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0735 ps=0.77 w=0.42 l=0.15
X13 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2b_2 VNB VPB VPWR VGND A_N X B
X0 VPWR a_212_413# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_297_47# a_27_413# a_212_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 X a_212_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.22895 ps=1.745 w=1 l=0.15
X3 X a_212_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.101875 ps=0.99 w=0.65 l=0.15
X4 a_212_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.07665 ps=0.785 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VPWR B a_212_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22895 pd=1.745 as=0.0609 ps=0.71 w=0.42 l=0.15
X7 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND a_212_413# X VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_4 VNB VPB VGND VPWR A2 B1 Y A1
X0 a_28_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 a_462_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2 Y B1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4 a_462_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5 a_28_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 a_462_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.104 ps=0.97 w=0.65 l=0.15
X7 Y B1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y A1 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X11 a_28_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.145 ps=1.29 w=1 l=0.15
X12 VPWR A2 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X14 VGND A2 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X15 a_28_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X16 VPWR A1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X17 a_28_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 VGND A2 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X19 VPWR A2 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.155 ps=1.31 w=1 l=0.15
X20 a_28_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X21 Y A1 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X22 a_462_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X23 VPWR A1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211o_4 VNB VPB VGND VPWR A2 A1 C1 X B1
X0 X a_79_204# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR A1 a_473_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 a_473_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.195 ps=1.39 w=1 l=0.15
X3 X a_79_204# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X4 VGND C1 a_79_204# VNB sky130_fd_pr__nfet_01v8 ad=0.108875 pd=0.985 as=0.104 ps=0.97 w=0.65 l=0.15
X5 a_79_204# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.092625 ps=0.935 w=0.65 l=0.15
X6 VPWR a_79_204# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14 ps=1.28 w=1 l=0.15
X7 a_473_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14 ps=1.28 w=1 l=0.15
X8 a_473_297# B1 a_727_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.16 ps=1.32 w=1 l=0.15
X9 X a_79_204# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X10 VGND B1 a_79_204# VNB sky130_fd_pr__nfet_01v8 ad=0.13975 pd=1.08 as=0.12675 ps=1.04 w=0.65 l=0.15
X11 a_79_204# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.108875 ps=0.985 w=0.65 l=0.15
X12 VGND a_79_204# X VNB sky130_fd_pr__nfet_01v8 ad=0.092625 pd=0.935 as=0.095875 ps=0.945 w=0.65 l=0.15
X13 a_1123_47# A1 a_79_204# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X14 a_555_297# B1 a_473_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.26 ps=2.52 w=1 l=0.15
X15 VPWR A2 a_473_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X16 VGND A2 a_1123_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.091 ps=0.93 w=0.65 l=0.15
X17 a_951_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.13975 ps=1.08 w=0.65 l=0.15
X18 VPWR a_79_204# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND a_79_204# X VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X20 a_79_204# A1 a_951_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X21 a_79_204# C1 a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X22 a_727_297# C1 a_79_204# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X23 X a_79_204# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2b_4 VNB VPB VGND VPWR Y B_N A
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_27_297# a_419_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND a_419_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VGND a_419_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 Y a_419_21# a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X11 Y a_419_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VGND B_N a_419_21# VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.182 ps=1.86 w=0.65 l=0.15
X13 Y a_419_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VPWR B_N a_419_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.27 ps=2.54 w=1 l=0.15
X15 a_27_297# a_419_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 Y a_419_21# a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4bb_1 VPWR VGND VPB VNB B A X D_N C_N
X0 VGND A a_311_413# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 VPWR A a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.05985 ps=0.705 w=0.42 l=0.15
X2 a_393_413# a_205_93# a_311_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1215 pd=1.33 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND C_N a_27_410# VNB sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VPWR C_N a_27_410# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1226 pd=1.32 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 X a_311_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X6 VGND a_27_410# a_311_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.05985 ps=0.705 w=0.42 l=0.15
X7 a_561_297# B a_489_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.05985 pd=0.705 as=0.0441 ps=0.63 w=0.42 l=0.15
X8 a_205_93# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06195 ps=0.715 w=0.42 l=0.15
X9 a_205_93# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.1226 ps=1.32 w=0.42 l=0.15
X10 a_489_297# a_27_410# a_393_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1215 ps=1.33 w=0.42 l=0.15
X11 a_311_413# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 a_311_413# a_205_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.05985 pd=0.705 as=0.1092 ps=1.36 w=0.42 l=0.15
X13 X a_311_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.101875 ps=0.99 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor4b_1 VPB VNB VGND VPWR D_N C Y B A
X0 Y a_91_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_91_199# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR A a_341_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X6 a_245_297# C a_161_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X7 a_341_297# B a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X8 a_91_199# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X9 a_161_297# a_91_199# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.52 ps=3.04 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221o_2 VPWR VGND VPB VNB C1 B2 B1 A1 A2 X
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X1 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1575 ps=1.315 w=1 l=0.15
X3 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.102375 ps=0.965 w=0.65 l=0.15
X6 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X7 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X8 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X9 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X10 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X13 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3b_2 VGND VPWR VNB VPB X C B A_N
X0 a_109_53# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 X a_215_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12715 ps=1.095 w=0.65 l=0.15
X2 a_109_53# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND C a_373_53# VNB sky130_fd_pr__nfet_01v8 ad=0.12715 pd=1.095 as=0.05355 ps=0.675 w=0.42 l=0.15
X4 VGND a_215_311# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR C a_215_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X6 VPWR a_215_311# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 X a_215_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X8 a_301_53# a_109_53# a_215_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_215_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_373_53# B a_301_53# VNB sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X11 VPWR a_109_53# a_215_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkinv_4 VNB VPB VPWR VGND A Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.1659 pd=1.63 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.14 ps=1.28 w=1 l=0.15
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.305 ps=2.61 w=1 l=0.15
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1386 ps=1.5 w=0.42 l=0.15
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o32a_1 VPB VNB VPWR VGND X A1 A2 A3 B2 B1
X0 a_77_199# B2 a_227_47# VNB sky130_fd_pr__nfet_01v8 ad=0.13325 pd=1.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X1 a_323_297# A2 a_227_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.165 ps=1.33 w=1 l=0.15
X2 a_227_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3 a_227_47# B1 a_77_199# VNB sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.13325 ps=1.06 w=0.65 l=0.15
X4 VGND a_77_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VPWR B1 a_539_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.205 ps=1.41 w=1 l=0.15
X6 a_227_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X7 VPWR a_77_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=2.67 w=1 l=0.15
X8 a_77_199# A3 a_323_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X9 VGND A2 a_227_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.10725 ps=0.98 w=0.65 l=0.15
X10 a_227_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_539_297# B2 a_77_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=1.41 as=0.195 ps=1.39 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_8 VPB VNB VGND VPWR A X
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X21 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221o_4 VNB VPB VPWR VGND A2 X A1 C1 B1 B2
X0 VGND A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VGND B2 a_1053_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_804_297# B1 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=1.69 as=0.135 ps=1.27 w=1 l=0.15
X3 a_79_21# A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_445_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_804_297# C1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_445_297# B1 a_804_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_1053_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_79_21# C1 a_804_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X10 a_1053_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_445_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 VGND C1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_804_297# B2 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X18 a_79_21# B1 a_1053_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_79_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_445_297# B2 a_804_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.345 ps=1.69 w=1 l=0.15
X21 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 a_445_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 a_445_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.135 ps=1.27 w=1 l=0.15
X24 VPWR A2 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 VPWR A1 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1375 ps=1.275 w=1 l=0.15
X26 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X27 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a41o_2 VNB VPB VGND VPWR X A1 A2 A3 A4 B1
X0 a_381_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR A2 a_381_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.215 ps=1.43 w=1 l=0.15
X2 a_465_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_549_47# A3 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.13975 pd=1.08 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_665_47# A2 a_549_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13975 ps=1.08 w=0.65 l=0.15
X7 a_381_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.215 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A4 a_381_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_381_297# B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 a_79_21# A1 a_665_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2_4 VNB VPB VGND VPWR A X B
X0 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X1 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VGND B a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 a_110_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X8 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X11 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22oi_1 VPWR VGND VPB VNB B2 B1 Y A1 A2
X0 Y B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X1 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.135 ps=1.27 w=1 l=0.15
X3 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 a_381_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_109_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X7 VGND A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.234 pd=2.02 as=0.06825 ps=0.86 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31a_2 VGND VPWR VPB VNB X A1 A2 A3 B1
X0 a_108_21# B1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X1 a_346_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 X a_108_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.26325 ps=2.11 w=0.65 l=0.15
X3 a_108_21# A3 a_430_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.425 as=0.165 ps=1.33 w=1 l=0.15
X4 a_430_297# A2 a_346_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR a_108_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.175 ps=1.35 w=1 l=0.15
X6 a_346_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND A2 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 X a_108_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.405 ps=2.81 w=1 l=0.15
X9 VPWR B1 a_108_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.2125 ps=1.425 w=1 l=0.15
X10 VGND a_108_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.11375 ps=1 w=0.65 l=0.15
X11 a_346_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12675 ps=1.04 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4b_1 VGND VPWR C A_N X D B VPB VNB
X0 a_297_47# a_27_47# a_193_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 a_369_47# B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 VPWR D a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.06615 ps=0.735 w=0.42 l=0.15
X3 X a_193_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1034 ps=1 w=0.65 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VGND D a_469_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1034 pd=1 as=0.0609 ps=0.71 w=0.42 l=0.15
X6 X a_193_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X7 VPWR B a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X8 a_193_413# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.1281 ps=1.03 w=0.42 l=0.15
X9 a_193_413# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_469_47# C a_369_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0735 ps=0.77 w=0.42 l=0.15
X11 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a311o_2 VPB VNB VGND VPWR C1 B1 A1 A2 A3 X
X0 a_79_21# C1 a_635_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.21 ps=1.42 w=1 l=0.15
X1 VPWR A2 a_319_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.17 ps=1.34 w=1 l=0.15
X2 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.13975 pd=1.08 as=0.13325 ps=1.06 w=0.65 l=0.15
X3 a_417_47# A2 a_319_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12025 pd=1.02 as=0.1105 ps=0.99 w=0.65 l=0.15
X4 a_79_21# A1 a_417_47# VNB sky130_fd_pr__nfet_01v8 ad=0.13325 pd=1.06 as=0.12025 ps=1.02 w=0.65 l=0.15
X5 a_319_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1105 pd=0.99 as=0.156 ps=1.13 w=0.65 l=0.15
X6 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.24 pd=1.48 as=0.135 ps=1.27 w=1 l=0.15
X7 a_319_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.185 ps=1.37 w=1 l=0.15
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.156 pd=1.13 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_319_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.34 as=0.24 ps=1.48 w=1 l=0.15
X10 a_79_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13975 ps=1.08 w=0.65 l=0.15
X11 a_635_297# B1 a_319_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.21 ps=1.42 w=1 l=0.15
X12 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2111oi_4 VNB VPB VGND VPWR A1 Y D1 C1 A2 B1
X0 Y D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_455_297# B1 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.26 ps=2.52 w=1 l=0.15
X2 a_28_297# D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 a_821_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4 a_28_297# C1 a_455_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 a_455_297# C1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.091 ps=0.93 w=0.65 l=0.15
X7 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 VPWR A2 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.2 ps=1.4 w=1 l=0.15
X9 Y D1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X10 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X11 VGND D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 Y D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X13 a_821_297# B1 a_455_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X15 Y D1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.117 ps=1.01 w=0.65 l=0.15
X17 a_1205_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X18 a_28_297# C1 a_455_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14 ps=1.28 w=1 l=0.15
X19 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.12675 ps=1.04 w=0.65 l=0.15
X20 a_1205_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X21 a_821_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.14 ps=1.28 w=1 l=0.15
X22 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X23 Y A1 a_1205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X24 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X25 VPWR A1 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.145 ps=1.29 w=1 l=0.15
X26 Y A1 a_1205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.182 ps=1.86 w=0.65 l=0.15
X27 a_1205_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.121875 pd=1.025 as=0.091 ps=0.93 w=0.65 l=0.15
X28 a_28_297# D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X29 VGND A2 a_1205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X30 a_455_297# B1 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X31 a_821_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2 pd=1.4 as=0.15 ps=1.3 w=1 l=0.15
X32 a_1205_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X33 VGND A2 a_1205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.121875 ps=1.025 w=0.65 l=0.15
X34 VPWR A1 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.14 ps=1.28 w=1 l=0.15
X35 a_821_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X36 VPWR A2 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X37 a_455_297# C1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X38 a_821_297# B1 a_455_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X39 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o221ai_1 VPB VNB VGND VPWR A1 A2 Y B2 C1 B1
X0 a_109_47# B1 a_213_123# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1652 ps=1.82 w=0.65 l=0.15
X1 Y B2 a_295_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.12 ps=1.24 w=1 l=0.15
X2 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3 a_213_123# B2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_295_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12 pd=1.24 as=0.38 ps=1.76 w=1 l=0.15
X5 a_493_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.225 ps=1.45 w=1 l=0.15
X6 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=1.76 as=0.28 ps=2.56 w=1 l=0.15
X7 VGND A2 a_213_123# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.117 ps=1.01 w=0.65 l=0.15
X8 a_213_123# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_109_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.1654 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ba_4 VNB VPB VGND VPWR B1_N X A2 A1
X0 VPWR B1_N a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.38 ps=2.76 w=1 l=0.15
X1 VPWR A1 a_743_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_743_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X3 a_575_47# a_27_297# a_187_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_743_297# A2 a_187_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR a_27_297# a_187_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6 a_187_21# A2 a_743_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 a_187_21# a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_187_21# a_27_297# a_575_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9 VGND B1_N a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.19825 ps=1.91 w=0.65 l=0.15
X10 VGND A2 a_575_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VPWR a_187_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VGND A1 a_575_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VGND a_187_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 X a_187_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VPWR a_187_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_575_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_575_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 X a_187_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 X a_187_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 X a_187_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 VGND a_187_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31ai_1 VPB VNB A1 A2 A3 Y B1 VPWR VGND
X0 Y B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.19825 ps=1.26 w=0.65 l=0.15
X1 Y A3 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3925 pd=1.785 as=0.135 ps=1.27 w=1 l=0.15
X2 a_193_297# A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.3925 ps=1.785 w=1 l=0.15
X5 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 a_109_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_2 VPWR VGND VPB VNB B D C A X
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.101875 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.91 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14825 ps=1.34 w=1 l=0.15
X9 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31oi_1 VGND VPWR VPB VNB A3 A2 A1 Y B1
X0 Y A1 a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.118625 ps=1.015 w=0.65 l=0.15
X1 a_181_47# A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.06825 ps=0.86 w=0.65 l=0.15
X2 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.105625 ps=0.975 w=0.65 l=0.15
X3 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.135 ps=1.27 w=1 l=0.15
X4 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1625 ps=1.325 w=1 l=0.15
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.1525 ps=1.305 w=1 l=0.15
X6 a_109_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3b_1 VPB VNB VGND VPWR C_N B Y A
X0 VGND a_91_199# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VPWR A a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X3 a_91_199# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_245_297# B a_161_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_91_199# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X7 a_161_297# a_91_199# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21a_2 VNB VPB VGND VPWR X B1 A2 A1
X0 VPWR A1 a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.16 ps=1.32 w=1 l=0.15
X1 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.4 ps=1.8 w=1 l=0.15
X2 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.089375 ps=0.925 w=0.65 l=0.15
X3 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X4 a_470_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.4 pd=1.8 as=0.1375 ps=1.275 w=1 l=0.15
X6 a_384_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X7 a_384_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.104 ps=0.97 w=0.65 l=0.15
X8 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X9 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2b_4 VNB VPB VGND VPWR X A B_N
X0 VPWR a_219_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND B_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0.201775 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VPWR A a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.34 as=0.105 ps=1.21 w=1 l=0.15
X3 a_27_53# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 X a_219_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1105 ps=0.99 w=0.65 l=0.15
X5 a_301_297# a_27_53# a_219_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X6 X a_219_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND A a_219_297# VNB sky130_fd_pr__nfet_01v8 ad=0.1105 pd=0.99 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR a_219_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND a_219_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 X a_219_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.17 ps=1.34 w=1 l=0.15
X11 VGND a_219_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.96 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_219_297# a_27_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.201775 ps=1.4 w=0.65 l=0.15
X13 X a_219_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3b_4 VNB VPB VGND VPWR B C A_N Y
X0 VGND C a_633_47# VNB sky130_fd_pr__nfet_01v8 ad=0.234 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_633_47# B a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_633_47# B a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 a_215_47# B a_633_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_215_47# B a_633_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_633_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X17 a_633_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X20 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X22 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X23 VGND C a_633_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X25 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor4_2 VNB VPB VGND VPWR B D Y A C
X0 a_281_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_475_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y D a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND D Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X9 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X12 a_475_297# C a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_281_297# C a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X14 a_27_297# B a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X15 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor4b_4 VPB VNB VGND VPWR B D_N A C Y
X0 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VGND D_N a_1191_21# VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_803_297# a_1191_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 a_445_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 Y a_1191_21# a_803_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_803_297# a_1191_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 Y a_1191_21# a_803_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25675 ps=1.44 w=0.65 l=0.15
X12 Y a_1191_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VPWR D_N a_1191_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_27_297# B a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X19 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 VGND a_1191_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 VGND a_1191_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 a_445_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 a_803_297# C a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X27 a_27_297# B a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 a_445_297# C a_803_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 a_803_297# C a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 Y a_1191_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X32 a_445_297# C a_803_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X33 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4bb_4 VNB VPB VGND VPWR A_N C D X B_N
X0 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X1 a_174_21# a_832_21# a_766_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_832_21# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1764 ps=1.68 w=0.42 l=0.15
X4 a_766_47# a_27_47# a_652_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.1365 ps=1.07 w=0.65 l=0.15
X5 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14075 ps=1.325 w=1 l=0.15
X7 VPWR B_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_652_47# C a_556_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.07 as=0.10725 ps=0.98 w=0.65 l=0.15
X9 a_832_21# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.31165 ps=2.125 w=0.42 l=0.15
X10 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X11 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_556_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.11375 ps=1 w=0.65 l=0.15
X13 a_174_21# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.175 ps=1.35 w=1 l=0.15
X14 VPWR C a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.165 ps=1.33 w=1 l=0.15
X15 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VPWR a_832_21# a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31165 pd=2.125 as=0.165 ps=1.33 w=1 l=0.15
X18 a_174_21# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.21 ps=1.42 w=1 l=0.15
X19 VGND B_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_8 VNB VPB VGND VPWR A Y B
X0 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.135 ps=1.27 w=1 l=0.15
X24 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X29 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X31 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21a_4 VNB VPB VPWR VGND A2 A1 X B1
X0 X a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_475_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2 X a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X4 a_762_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.31 ps=1.62 w=1 l=0.15
X5 a_475_47# B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.091 ps=0.93 w=0.65 l=0.15
X6 VGND A2 a_475_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X7 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 X a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X10 a_80_21# A2 a_762_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_80_21# B1 a_475_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X12 a_80_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15 ps=1.3 w=1 l=0.15
X13 a_475_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.117 ps=1.01 w=0.65 l=0.15
X14 X a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 VPWR A1 a_934_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X16 a_934_297# A2 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X17 VPWR B1 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=1.62 as=0.14 ps=1.28 w=1 l=0.15
X18 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND A1 a_475_47# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.117 ps=1.01 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3b_2 VNB VPB VGND VPWR A_N C B Y
X0 a_408_47# B a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_408_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y a_27_47# a_408_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17575 pd=1.395 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VGND C a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6 a_218_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11975 ps=1.045 w=0.65 l=0.15
X7 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 a_218_47# B a_408_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.17575 ps=1.395 w=1 l=0.15
X12 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11975 pd=1.045 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211oi_2 VPWR VGND VPB VNB A2 A1 Y B1 C1
X0 VGND A2 a_485_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1 VPWR A1 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 a_37_297# B1 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4 a_485_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X5 a_292_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X7 VPWR A2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8 a_485_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X11 a_37_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 Y A1 a_485_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X13 Y C1 a_37_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X14 a_292_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X15 a_292_297# B1 a_37_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor4_1 VPB VNB VGND VPWR Y D C B A
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.089375 ps=0.925 w=0.65 l=0.15
X1 a_191_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.13 ps=1.26 w=1 l=0.15
X2 VPWR A a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.118625 ps=1.015 w=0.65 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_297_297# B a_191_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X6 a_109_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.26 as=0.26 ps=2.52 w=1 l=0.15
X7 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a311oi_1 VPB VNB Y C1 B1 A1 A2 A3 VPWR VGND
X0 Y A1 a_194_47# VNB sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_194_47# A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X2 Y C1 a_376_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1725 ps=1.345 w=1 l=0.15
X3 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X4 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.112125 ps=0.995 w=0.65 l=0.15
X5 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.115375 ps=1.005 w=0.65 l=0.15
X6 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X7 a_376_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.165 ps=1.33 w=1 l=0.15
X8 a_109_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X9 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3b_2 VPB VNB VGND VPWR A Y C_N B
X0 a_281_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND a_531_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR C_N a_531_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X7 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X9 a_281_297# a_531_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X10 Y a_531_21# a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X11 VGND C_N a_531_21# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X12 a_27_297# B a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X13 Y a_531_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand4_1 VPB VNB VPWR VGND A C D Y B
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X2 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_47# C a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y A a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X5 a_277_47# B a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 a_109_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt tt_um_MichaelBell_tinyQV VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2]
+ ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3]
+ uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3]
+ uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3]
+ uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3]
+ uo_out[4] uo_out[5] uo_out[6] uo_out[7]
XFILLER_0_27_82 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7963_ i_tinyqv.cpu.i_core.mepc\[23\] clknet_leaf_35_clk _0100_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_6914_ VPWR VGND VGND VPWR _3260_ _3268_ net16 sky130_fd_sc_hd__nor2_2
X_7894_ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[17\] clknet_leaf_2_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[17\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6845_ VPWR VGND VGND VPWR _3216_ i_tinyqv.cpu.instr_data_start\[21\] i_tinyqv.cpu.imm\[21\]
+ sky130_fd_sc_hd__or2_1
X_6776_ VPWR VGND VGND VPWR _0881_ _3153_ i_tinyqv.cpu.imm\[15\] sky130_fd_sc_hd__nand2_1
X_3988_ VPWR VGND _0839_ _0614_ i_tinyqv.cpu.counter\[4\] VPWR VGND sky130_fd_sc_hd__and2_1
X_5727_ VGND VPWR _2374_ _2372_ _2181_ _2373_ VPWR VGND sky130_fd_sc_hd__and3_1
X_8515_ i_tinyqv.cpu.i_core.i_instrret.register\[21\] clknet_leaf_45_clk i_tinyqv.cpu.i_core.i_instrret.reg_buf\[21\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_8446_ i_tinyqv.cpu.imm\[24\] clknet_leaf_8_clk _0544_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5658_ VGND VPWR _0168_ _2323_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5589_ VGND VPWR VPWR VGND i_uart_rx.cycle_counter\[10\] i_uart_rx.cycle_counter\[8\]
+ i_uart_rx.cycle_counter\[9\] _2273_ sky130_fd_sc_hd__or3b_1
X_8377_ i_debug_uart_tx.uart_tx_data\[2\] clknet_leaf_25_clk _0475_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_4609_ VPWR VGND VGND VPWR _1445_ i_tinyqv.cpu.instr_data\[3\]\[3\] _1422_ sky130_fd_sc_hd__or2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.i_regbuf\[25\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[25\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[29\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7328_ VPWR VGND VPWR VGND _0711_ i_tinyqv.cpu.mem_op_increment_reg _0660_ _3596_
+ sky130_fd_sc_hd__a21oi_1
X_7259_ VPWR VGND VGND VPWR _3334_ _3539_ _3301_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_51_556 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xrebuffer7 VPWR VGND VPWR VGND net323 _0651_ sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_51_578 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_51_567 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_4960_ VPWR VGND VPWR VGND _1727_ net238 _1735_ _0004_ sky130_fd_sc_hd__a21o_1
X_4891_ VGND VPWR VPWR VGND _1689_ _1638_ _1685_ net152 sky130_fd_sc_hd__mux2_1
X_3911_ VGND VPWR VPWR VGND _0654_ _0762_ _0754_ _0763_ sky130_fd_sc_hd__mux2_2
X_6630_ VGND VPWR VPWR VGND _3021_ _3023_ _3022_ sky130_fd_sc_hd__xor2_1
X_3842_ VGND VPWR _0694_ _0608_ _0614_ i_tinyqv.cpu.imm\[31\] VPWR VGND sky130_fd_sc_hd__and3_1
X_6561_ VGND VPWR VGND VPWR _2969_ _2966_ _2968_ _2929_ _2956_ sky130_fd_sc_hd__a211o_1
XFILLER_0_27_542 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_5512_ VGND VPWR _2218_ _2200_ _2220_ net102 VPWR VGND sky130_fd_sc_hd__o21ai_1
X_8300_ i_tinyqv.mem.q_ctrl.is_writing clknet_leaf_16_clk _0399_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_95 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_3773_ VPWR VGND _0625_ i_tinyqv.cpu.i_core.i_registers.rs1\[2\] VPWR VGND sky130_fd_sc_hd__buf_6
X_6492_ VPWR VGND VGND VPWR i_tinyqv.mem.q_ctrl.data_req _2906_ _0868_ sky130_fd_sc_hd__nand2_4
XFILLER_0_14_247 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5443_ VGND VPWR VGND VPWR _1725_ _0997_ _2169_ _0991_ sky130_fd_sc_hd__nand3_4
XFILLER_0_14_269 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_42_589 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_8231_ i_tinyqv.cpu.i_core.mepc\[2\] clknet_leaf_34_clk _0331_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_2
X_8162_ i_tinyqv.cpu.instr_data\[2\]\[11\] clknet_leaf_11_clk _0274_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5374_ VGND VPWR _2106_ _2107_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_4325_ VPWR VGND VGND VPWR _1171_ _1172_ _0745_ sky130_fd_sc_hd__nand2_1
X_7113_ VGND VPWR VGND VPWR _3421_ _3416_ _3419_ _1460_ _3420_ sky130_fd_sc_hd__a211o_1
X_8093_ gpio_out\[4\] clknet_leaf_18_clk _0004_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_464 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4256_ VGND VPWR i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt\[0\] _1103_ VPWR
+ VGND sky130_fd_sc_hd__clkbuf_4
X_7044_ VGND VPWR VGND VPWR _0519_ net209 _3282_ _3357_ _1753_ sky130_fd_sc_hd__o211a_1
X_4187_ VPWR VGND VGND VPWR _1033_ _0877_ _1034_ sky130_fd_sc_hd__nor2_1
X_7946_ i_tinyqv.cpu.i_core.load_done clknet_leaf_51_clk net139 VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_7877_ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[0\] clknet_leaf_48_clk _0062_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6828_ VPWR VGND VGND VPWR _3040_ _3201_ _3051_ _3200_ _3199_ sky130_fd_sc_hd__o211ai_1
X_6759_ VPWR VGND VGND VPWR _3136_ _3138_ _3137_ sky130_fd_sc_hd__nand2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.i_regbuf\[26\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[26\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[30\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_8429_ i_tinyqv.cpu.i_core.imm_lo\[7\] clknet_leaf_22_clk _0527_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_33_567 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold170 net199 i_uart_rx.cycle_counter\[7\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 net210 i_tinyqv.mem.q_ctrl.spi_ram_b_select VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 net221 i_tinyqv.cpu.i_core.imm_lo\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_55_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.i_regbuf\[25\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[25\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[29\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_cycles.i_regbuf\[23\] i_tinyqv.cpu.i_core.i_cycles.reg_buf\[23\]
+ i_tinyqv.cpu.i_core.i_cycles.register\[27\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4110_ VGND VPWR _0865_ _0957_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_5090_ VGND VPWR _1849_ _1850_ _1847_ VPWR VGND sky130_fd_sc_hd__xnor2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.i_regbuf\[14\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[14\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[18\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4041_ VGND VPWR VGND VPWR _0885_ i_tinyqv.cpu.instr_len\[1\] _0749_ _0887_ _0888_
+ sky130_fd_sc_hd__a31o_2
X_7800_ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[19\] clknet_leaf_0_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[19\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5992_ VGND VPWR _0264_ _2560_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4943_ VPWR VGND _1724_ net1 i_tinyqv.mem.q_ctrl.spi_data_oe\[0\] VPWR VGND sky130_fd_sc_hd__and2_1
X_7731_ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[14\] clknet_leaf_0_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[14\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7662_ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[9\] clknet_leaf_55_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[9\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6613_ VGND VPWR _3008_ _3009_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_4874_ VGND VPWR VGND VPWR i_tinyqv.cpu.i_core.i_registers.rd\[2\] i_tinyqv.cpu.i_core.i_registers.rd\[1\]
+ _1679_ i_tinyqv.cpu.i_core.i_registers.rd\[0\] sky130_fd_sc_hd__nand3_2
XFILLER_0_61_117 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7593_ i_tinyqv.cpu.i_core.i_registers.reg_access\[13\]\[0\] clknet_leaf_1_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[4\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_3825_ VGND VPWR VGND VPWR _0677_ i_tinyqv.cpu.i_core.i_registers.rs2\[3\] i_tinyqv.cpu.i_core.i_registers.rs2\[2\]
+ net37 net38 sky130_fd_sc_hd__and4_2
X_6544_ VPWR VGND VGND VPWR _2954_ i_debug_uart_tx.uart_tx_data\[4\] _2909_ sky130_fd_sc_hd__or2_1
X_3756_ VGND VPWR i_tinyqv.cpu.counter\[2\] _0608_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_266 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6475_ VPWR VGND _2897_ _2896_ VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_0_15_556 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_40_93 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_71_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_8214_ i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt\[1\] clknet_leaf_39_clk _0326_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_5426_ VPWR VGND _2155_ _1448_ VPWR VGND sky130_fd_sc_hd__buf_2
X_8145_ i_tinyqv.cpu.data_addr\[20\] clknet_leaf_32_clk _0257_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_5357_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.mepc\[1\] net18 _2093_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_58_Left_139 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5288_ VGND VPWR _2014_ _2011_ _2040_ _2013_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_8076_ debug_rd_r\[0\] clknet_leaf_51_clk i_tinyqv.cpu.debug_rd\[0\] VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_4308_ VGND VPWR VPWR VGND _1155_ _1064_ _1103_ _1062_ sky130_fd_sc_hd__mux2_1
X_4239_ VGND VPWR VPWR VGND _1086_ i_tinyqv.cpu.i_core.i_shift.a\[31\] _1036_ i_tinyqv.cpu.i_core.i_shift.a\[0\]
+ sky130_fd_sc_hd__mux2_1
X_7027_ VGND VPWR _3343_ _3281_ _3341_ _3342_ VPWR VGND sky130_fd_sc_hd__and3_1
X_7929_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[20\] clknet_leaf_36_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[20\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_67_Left_148 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_80_415 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_45_180 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_61_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_33_364 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_76_Left_157 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.i_regbuf\[30\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[30\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[2\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_309 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4590_ VGND VPWR VPWR VGND _1426_ _1425_ _1416_ _1421_ _1423_ sky130_fd_sc_hd__a31oi_4
X_6260_ VPWR VGND VPWR VGND _2734_ _0872_ _2735_ _2736_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5211_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[11\] _1966_ _1845_ sky130_fd_sc_hd__nand2_1
X_6191_ VGND VPWR _0347_ _2676_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5142_ VPWR VGND VGND VPWR _1871_ _1900_ _1874_ sky130_fd_sc_hd__nand2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.i_regbuf\[15\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[15\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[19\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5073_ VPWR VGND VPWR VGND _1789_ i_tinyqv.cpu.i_core.i_shift.a\[5\] _1309_ _1833_
+ i_tinyqv.cpu.i_core.i_shift.a\[4\] sky130_fd_sc_hd__a22o_1
X_4024_ VGND VPWR _0082_ _0873_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5975_ VGND VPWR VPWR VGND _2549_ _2548_ _2501_ i_tinyqv.cpu.data_addr\[22\] sky130_fd_sc_hd__mux2_1
X_4926_ VPWR VGND _1711_ _1710_ VPWR VGND sky130_fd_sc_hd__buf_2
X_7714_ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[29\] clknet_leaf_56_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[29\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4857_ VGND VPWR VPWR VGND _1670_ i_tinyqv.cpu.debug_rd\[0\] _1669_ i_tinyqv.cpu.i_core.i_registers.reg_access\[9\]\[0\]
+ sky130_fd_sc_hd__mux2_1
X_7645_ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[24\] clknet_leaf_57_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[24\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7576_ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[19\] clknet_leaf_58_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[19\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_3808_ VPWR VGND _0660_ i_tinyqv.cpu.i_core.i_registers.rs2\[2\] VPWR VGND sky130_fd_sc_hd__buf_2
X_6527_ VGND VPWR VPWR VGND _2939_ _2938_ _2916_ net12 sky130_fd_sc_hd__mux2_1
X_4788_ VGND VPWR VPWR VGND _1623_ _1622_ _0908_ _1621_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_364 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6458_ VGND VPWR _0407_ _2883_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xi_tinyqv.cpu.i_core.i_instrret.i_regbuf\[9\] i_tinyqv.cpu.i_core.i_instrret.reg_buf\[9\]
+ i_tinyqv.cpu.i_core.i_instrret.register\[13\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6389_ VGND VPWR _2823_ _2787_ _2828_ _2804_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_5409_ VPWR VGND VGND VPWR _2134_ _2138_ _2139_ sky130_fd_sc_hd__nor2_1
X_8128_ i_tinyqv.cpu.data_addr\[3\] clknet_leaf_28_clk _0240_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_592 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_8059_ i_spi.bits_remaining\[1\] clknet_leaf_28_clk _0194_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_570 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5760_ VGND VPWR _0192_ _2401_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5691_ VGND VPWR VGND VPWR _0176_ i_debug_uart_tx.uart_tx_data\[3\] _2330_ _2348_
+ _2299_ sky130_fd_sc_hd__o211a_1
X_4711_ VGND VPWR VGND VPWR _1480_ _1188_ net6 _1399_ _1546_ net5 _1547_ sky130_fd_sc_hd__mux4_1
X_7430_ VPWR VGND VPWR VGND _3632_ _3141_ _3678_ _3675_ _3677_ _2877_ sky130_fd_sc_hd__a221o_1
X_4642_ VPWR VGND VGND VPWR _1477_ _1478_ _1469_ sky130_fd_sc_hd__nor2_2
X_4573_ VPWR VGND _1409_ _1408_ VPWR VGND sky130_fd_sc_hd__buf_4
X_7361_ VPWR VGND VPWR VGND _3620_ _3618_ _2067_ _0573_ sky130_fd_sc_hd__a21oi_1
X_6312_ VGND VPWR _0378_ _2766_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7292_ VPWR VGND _3567_ _3564_ _2124_ _3291_ _3566_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_6243_ VPWR VGND VGND VPWR _2704_ _2721_ _2722_ sky130_fd_sc_hd__nor2_1
X_6174_ VGND VPWR VPWR VGND _2668_ i_tinyqv.cpu.i_core.mepc\[14\] _2667_ i_tinyqv.cpu.i_core.mepc\[10\]
+ sky130_fd_sc_hd__mux2_1
X_5125_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[9\] _1883_ _1167_ sky130_fd_sc_hd__nand2_1
X_5056_ VGND VPWR _1816_ _1817_ i_tinyqv.cpu.i_core.multiplier.accum\[6\] VPWR VGND
+ sky130_fd_sc_hd__xnor2_1
X_4007_ VGND VPWR VPWR VGND i_tinyqv.cpu.debug_instr_valid _0858_ i_tinyqv.cpu.is_jal
+ i_tinyqv.cpu.is_jalr sky130_fd_sc_hd__o21ai_4
X_5958_ VGND VPWR _0253_ _2537_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4909_ VGND VPWR _0060_ _1699_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5889_ VGND VPWR VPWR VGND _2490_ i_spi.data\[2\] _2386_ i_debug_uart_tx.uart_tx_data\[3\]
+ sky130_fd_sc_hd__mux2_1
X_7628_ i_tinyqv.cpu.i_core.i_registers.reg_access\[12\]\[3\] clknet_leaf_44_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[7\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.i_regbuf\[5\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[5\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[9\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7559_ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[2\] clknet_leaf_47_clk _0052_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_120 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.i_regbuf\[15\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[15\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[19\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 net103 i_tinyqv.cpu.i_core.i_registers.reg_access\[12\]\[2\] VPWR VGND VGND
+ VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 net92 i_tinyqv.cpu.i_core.i_instrret.data\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold96 net125 i_tinyqv.cpu.data_out\[15\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 net114 i_tinyqv.cpu.data_out\[28\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_448 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XANTENNA_5 _1729_ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xrebuffer17 VGND VPWR net46 _0643_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6930_ VPWR VGND VPWR VGND _3272_ _3253_ _3267_ _0490_ net140 sky130_fd_sc_hd__a22o_1
Xrebuffer28 VGND VPWR net57 _0645_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xrebuffer39 VGND VPWR net68 _0762_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6861_ VPWR VGND VGND VPWR _3231_ _3028_ _3230_ sky130_fd_sc_hd__or2_1
X_6792_ VPWR VGND VGND VPWR _3166_ _3168_ _3167_ sky130_fd_sc_hd__nand2_1
X_5812_ VPWR VGND VPWR VGND _0205_ _2083_ _2440_ _2431_ _2436_ sky130_fd_sc_hd__a211oi_1
X_5743_ VPWR VGND VGND VPWR _2387_ _2386_ i_spi.clock_count\[0\] sky130_fd_sc_hd__or2_1
X_8531_ i_tinyqv.cpu.i_core.cycle_count\[0\] clknet_leaf_50_clk i_tinyqv.cpu.i_core.i_cycles.reg_buf\[4\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5674_ VPWR VGND VPWR VGND _2335_ _2334_ sky130_fd_sc_hd__inv_2
X_8462_ i_tinyqv.cpu.i_core.i_registers.rs1\[1\] clknet_leaf_51_clk _0560_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_8393_ i_tinyqv.cpu.data_out\[18\] clknet_leaf_26_clk _0491_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_7413_ _3664_ _2877_ _3660_ _3663_ _3004_ VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_4625_ VPWR VGND _1461_ _1416_ VPWR VGND sky130_fd_sc_hd__buf_4
X_7344_ VGND VPWR VPWR VGND _3608_ _2152_ i_tinyqv.cpu.additional_mem_ops\[0\] _2147_
+ sky130_fd_sc_hd__mux2_1
X_4556_ VPWR VGND VGND VPWR _1173_ _1392_ _0855_ sky130_fd_sc_hd__nor2_2
XFILLER_0_13_676 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_40_462 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7275_ VPWR VGND VGND VPWR net243 _3474_ _3552_ _0555_ sky130_fd_sc_hd__o21a_1
X_4487_ VPWR VGND VGND VPWR _1324_ _1326_ _1325_ sky130_fd_sc_hd__nand2_1
X_6226_ VPWR VGND _2706_ _2705_ _2704_ VPWR VGND sky130_fd_sc_hd__and2_1
X_6157_ VGND VPWR VPWR VGND _2659_ i_tinyqv.cpu.i_core.mepc\[6\] _2656_ i_tinyqv.cpu.i_core.mepc\[2\]
+ sky130_fd_sc_hd__mux2_1
X_5108_ VPWR VGND VGND VPWR _1054_ _1867_ _1845_ sky130_fd_sc_hd__nand2_1
X_6088_ VGND VPWR VPWR VGND _2612_ i_tinyqv.cpu.i_core.i_shift.a\[16\] _2596_ i_tinyqv.cpu.i_core.i_shift.a\[20\]
+ sky130_fd_sc_hd__mux2_1
X_5039_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[4\] _1801_ _1250_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_4410_ VGND VPWR VPWR VGND _0779_ _1178_ _0763_ _1253_ sky130_fd_sc_hd__or3b_1
X_5390_ VPWR VGND VGND VPWR _1483_ _2119_ _2120_ sky130_fd_sc_hd__nor2_1
X_4341_ VGND VPWR _1187_ _0846_ _0842_ _1025_ VPWR VGND sky130_fd_sc_hd__and3_1
X_4272_ VGND VPWR VGND VPWR _1048_ _1118_ _1077_ _1090_ _1100_ _1119_ sky130_fd_sc_hd__a311o_1
X_7060_ VPWR VGND VPWR VGND i_tinyqv.cpu.instr_data\[3\]\[4\] _3369_ _3373_ _3370_
+ i_tinyqv.cpu.instr_data\[2\]\[4\] _3372_ sky130_fd_sc_hd__a221o_1
X_6011_ VGND VPWR _0272_ _2571_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7962_ i_tinyqv.cpu.i_core.mepc\[22\] clknet_leaf_35_clk _0099_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_6913_ VGND VPWR VPWR VGND _0478_ _3267_ _3265_ _1619_ _3266_ net313 sky130_fd_sc_hd__a32o_1
X_7893_ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[16\] clknet_leaf_49_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[16\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6844_ VPWR VGND VGND VPWR i_tinyqv.cpu.instr_data_start\[21\] _3215_ i_tinyqv.cpu.imm\[21\]
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_359 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6775_ VPWR VGND VGND VPWR _3145_ _3152_ _3037_ i_tinyqv.cpu.instr_data_start\[14\]
+ _0455_ _1753_ sky130_fd_sc_hd__o221a_1
X_3987_ _0838_ _0608_ VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5726_ VPWR VGND VPWR VGND _2333_ i_debug_uart_tx.fsm_state\[0\] i_debug_uart_tx.fsm_state\[1\]
+ _2373_ sky130_fd_sc_hd__a21o_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.i_regbuf\[29\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[29\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[1\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_8514_ i_tinyqv.cpu.i_core.i_instrret.register\[20\] clknet_leaf_49_clk i_tinyqv.cpu.i_core.i_instrret.reg_buf\[20\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_8445_ i_tinyqv.cpu.imm\[23\] clknet_leaf_7_clk _0543_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_5657_ VGND VPWR VPWR VGND _2323_ _2322_ _2308_ i_tinyqv.cpu.instr_data\[3\]\[11\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_248 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5588_ VGND VPWR VGND VPWR _0149_ net191 _2263_ _2272_ _2240_ sky130_fd_sc_hd__o211a_1
X_8376_ i_debug_uart_tx.uart_tx_data\[1\] clknet_leaf_25_clk _0474_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_4608_ VPWR VGND VPWR VGND _1405_ _1438_ _1400_ _1444_ _1443_ sky130_fd_sc_hd__or4b_1
X_4539_ VGND VPWR VGND VPWR _1023_ _1022_ _1377_ _1378_ sky130_fd_sc_hd__o21ba_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.i_regbuf\[18\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[18\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[22\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7327_ VGND VPWR _3595_ i_tinyqv.cpu.mem_op_increment_reg _0660_ _0711_ VPWR VGND
+ sky130_fd_sc_hd__and3_1
X_7258_ VGND VPWR _0552_ _3538_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6209_ VGND VPWR _0351_ _2690_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7189_ VPWR VGND VPWR VGND _3438_ net227 _3486_ _0535_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_635 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xclkbuf_3_6__f_clk VGND VPWR VGND VPWR clknet_0_clk clknet_3_6__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_23_19 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_392 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xrebuffer8 VPWR VGND net37 i_tinyqv.cpu.i_core.i_registers.rs2\[1\] VPWR VGND sky130_fd_sc_hd__buf_6
X_3910_ VPWR VGND VGND VPWR _0761_ _0762_ _0757_ sky130_fd_sc_hd__nor2_2
X_4890_ VGND VPWR _0068_ _1688_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_104 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_3841_ VPWR VGND VPWR VGND i_tinyqv.cpu.i_core.imm_lo\[3\] _0689_ _0693_ _0691_ i_tinyqv.cpu.i_core.imm_lo\[11\]
+ _0692_ sky130_fd_sc_hd__a221o_1
XFILLER_0_39_370 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_6560_ VGND VPWR VGND VPWR _2968_ i_tinyqv.cpu.data_out\[22\] _2909_ _2914_ _2967_
+ sky130_fd_sc_hd__o211a_1
X_3772_ VPWR VGND _0624_ i_tinyqv.cpu.i_core.i_registers.rs1\[1\] VPWR VGND sky130_fd_sc_hd__buf_4
X_5511_ VPWR VGND VGND VPWR _2218_ net171 _0125_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_587 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6491_ VGND VPWR _0418_ _2905_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5442_ VGND VPWR VGND VPWR _0107_ _2153_ net252 _2168_ sky130_fd_sc_hd__a21bo_1
X_8230_ i_tinyqv.cpu.i_core.mepc\[1\] clknet_leaf_35_clk _0330_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_8161_ i_tinyqv.cpu.instr_data\[2\]\[10\] clknet_leaf_3_clk _0273_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5373_ VGND VPWR _2105_ _2106_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_8092_ gpio_out\[3\] clknet_leaf_18_clk _0003_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4324_ _1171_ _0746_ _0743_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_7112_ VPWR VGND VGND VPWR _3420_ _3299_ _3399_ _3350_ _3349_ _3292_ sky130_fd_sc_hd__o41a_1
X_7043_ VPWR VGND VGND VPWR _1495_ _3357_ _3282_ _3356_ _3342_ sky130_fd_sc_hd__o211ai_1
X_4255_ VGND VPWR VPWR VGND _1102_ i_tinyqv.cpu.i_core.i_shift.a\[9\] _1028_ i_tinyqv.cpu.i_core.i_shift.a\[22\]
+ sky130_fd_sc_hd__mux2_1
X_4186_ VPWR VGND VGND VPWR _1026_ _1032_ _1033_ sky130_fd_sc_hd__nor2_1
X_7945_ i_tinyqv.cpu.i_core.cy clknet_leaf_50_clk i_tinyqv.cpu.i_core.cy_out VPWR
+ VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7876_ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[31\] clknet_leaf_47_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[31\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6827_ VPWR VGND VGND VPWR _3040_ _3200_ _2542_ sky130_fd_sc_hd__nand2_1
X_6758_ VPWR VGND VGND VPWR _3137_ i_tinyqv.cpu.instr_data_start\[13\] i_tinyqv.cpu.imm\[13\]
+ sky130_fd_sc_hd__or2_1
X_5709_ _2360_ i_debug_uart_tx.cycle_counter\[0\] i_debug_uart_tx.cycle_counter\[2\]
+ i_debug_uart_tx.cycle_counter\[1\] _0989_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
X_6689_ VPWR VGND VGND VPWR _3051_ _3073_ _3074_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_481 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_8428_ i_tinyqv.cpu.i_core.imm_lo\[6\] clknet_leaf_9_clk _0526_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_2
X_8359_ i_tinyqv.cpu.instr_data_start\[17\] clknet_leaf_36_clk _0458_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.i_regbuf\[19\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[19\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[23\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold160 net189 i_tinyqv.mem.q_ctrl.addr\[18\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 net200 i_tinyqv.cpu.i_core.mie\[19\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 net211 i_tinyqv.cpu.i_core.mepc\[23\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 net222 i_tinyqv.cpu.i_core.mepc\[21\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.i_regbuf\[22\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[22\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[26\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_159 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_51_387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.i_regbuf\[18\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[18\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[22\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_cycles.i_regbuf\[16\] i_tinyqv.cpu.i_core.i_cycles.reg_buf\[16\]
+ i_tinyqv.cpu.i_core.i_cycles.register\[20\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4040_ VPWR VGND VGND VPWR _0887_ _0886_ _0885_ sky130_fd_sc_hd__nor2_4
X_5991_ VPWR VGND _2560_ _2559_ _2079_ VPWR VGND sky130_fd_sc_hd__and2_1
X_4942_ VGND VPWR _1723_ uio_out[5] VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_7730_ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[13\] clknet_leaf_54_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[13\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7661_ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[8\] clknet_leaf_0_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[8\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6612_ VPWR VGND VGND VPWR _3004_ _3007_ _3008_ sky130_fd_sc_hd__nor2_1
X_4873_ VGND VPWR _0077_ _1678_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7592_ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[3\] clknet_leaf_57_clk _0049_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_3824_ VPWR VGND VPWR VGND _0675_ i_tinyqv.cpu.i_core.i_registers.reg_access\[12\]\[3\]
+ _0674_ _0676_ i_tinyqv.cpu.i_core.i_registers.reg_access\[5\]\[3\] sky130_fd_sc_hd__a22o_1
X_6543_ VGND VPWR VPWR VGND _2953_ i_tinyqv.cpu.data_out\[20\] _2912_ i_tinyqv.cpu.data_out\[28\]
+ sky130_fd_sc_hd__mux2_1
X_3755_ VPWR VGND VPWR VGND _0607_ i_tinyqv.cpu.counter\[4\] sky130_fd_sc_hd__inv_2
XFILLER_0_15_546 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6474_ VPWR VGND VPWR VGND i_tinyqv.mem.q_ctrl.read_cycles_count\[0\] _2787_ _1713_
+ _2896_ _2782_ sky130_fd_sc_hd__or4b_1
XFILLER_0_42_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Right_12 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5425_ VGND VPWR _0104_ _2154_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8213_ i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt\[0\] clknet_leaf_40_clk _0325_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_2_473 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_8144_ i_tinyqv.cpu.data_addr\[19\] clknet_leaf_34_clk _0256_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_5356_ VPWR VGND VPWR VGND _2087_ net244 _0840_ _0097_ _2092_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5287_ VGND VPWR VPWR VGND _2037_ _2039_ _2038_ sky130_fd_sc_hd__xor2_1
X_4307_ VGND VPWR VPWR VGND _1154_ _1061_ _1103_ _1114_ sky130_fd_sc_hd__mux2_1
X_8075_ i_tinyqv.cpu.i_core.mie\[16\] clknet_leaf_37_clk _0210_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_4238_ VGND VPWR VPWR VGND _1085_ i_tinyqv.cpu.i_core.i_shift.a\[30\] _1036_ i_tinyqv.cpu.i_core.i_shift.a\[1\]
+ sky130_fd_sc_hd__mux2_1
X_7026_ VPWR VGND VPWR VGND _3287_ _3307_ _1514_ _3342_ sky130_fd_sc_hd__or3_1
X_4169_ VGND VPWR _1016_ i_tinyqv.cpu.data_write_n\[0\] i_tinyqv.cpu.data_read_n\[0\]
+ _1015_ VPWR VGND sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_21_Right_21 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7928_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[19\] clknet_leaf_36_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[19\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7859_ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[14\] clknet_leaf_2_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[14\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_30_Right_30 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_60_184 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_45_28 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.i_regbuf\[23\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[23\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[27\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_365 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_10_97 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5210_ VPWR VGND VGND VPWR _1963_ _1965_ _1964_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_560 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_6190_ VGND VPWR VPWR VGND _2676_ i_tinyqv.cpu.i_core.mepc\[22\] _2667_ i_tinyqv.cpu.i_core.mepc\[18\]
+ sky130_fd_sc_hd__mux2_1
X_5141_ VPWR VGND _1899_ _1898_ _1897_ VPWR VGND sky130_fd_sc_hd__and2_1
X_5072_ VPWR VGND VGND VPWR _1832_ _1807_ _1831_ sky130_fd_sc_hd__or2_1
X_4023_ VPWR VGND _0873_ _0872_ i_tinyqv.mem.q_ctrl.data_req VPWR VGND sky130_fd_sc_hd__and2_1
X_7713_ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[28\] clknet_leaf_0_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[28\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5974_ VGND VPWR VPWR VGND _2548_ i_tinyqv.cpu.i_core.mepc\[22\] _2106_ i_tinyqv.cpu.i_core.i_shift.a\[26\]
+ sky130_fd_sc_hd__mux2_1
X_4925_ i_tinyqv.mem.q_ctrl.fsm_state\[1\] i_tinyqv.mem.q_ctrl.fsm_state\[0\] _1710_
+ i_tinyqv.mem.q_ctrl.fsm_state\[2\] VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
XFILLER_0_74_243 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_7644_ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[23\] clknet_leaf_46_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[23\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4856_ VPWR VGND _1647_ _1669_ _1658_ VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_0_62_449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.i_regbuf\[11\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[11\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[15\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7575_ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[18\] clknet_leaf_54_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[18\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_3807_ VPWR VGND VPWR VGND net37 i_tinyqv.cpu.i_core.i_registers.rs2\[3\] net38 _0659_
+ i_tinyqv.cpu.i_core.i_registers.rs2\[2\] sky130_fd_sc_hd__or4b_1
X_6526_ VGND VPWR VPWR VGND _2938_ _2937_ _2914_ _2936_ sky130_fd_sc_hd__mux2_1
X_4787_ VGND VPWR VPWR VGND _1622_ i_tinyqv.mem.qspi_data_buf\[11\] _1017_ i_tinyqv.cpu.instr_data_in\[11\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_376 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_6457_ VPWR VGND _2883_ _2882_ _2832_ VPWR VGND sky130_fd_sc_hd__and2_1
X_6388_ VPWR VGND VPWR VGND _2824_ _2800_ _2826_ _2827_ sky130_fd_sc_hd__a21oi_1
X_5408_ VPWR VGND VGND VPWR _1490_ _2138_ _2128_ sky130_fd_sc_hd__nand2_1
X_8127_ i_tinyqv.cpu.data_addr\[2\] clknet_leaf_25_clk _0239_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_2
X_5339_ VGND VPWR _1752_ _2079_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_8058_ i_spi.bits_remaining\[0\] clknet_leaf_28_clk _0193_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7009_ VGND VPWR VGND VPWR _0514_ _3312_ _3325_ _3327_ _3205_ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_298 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_25_129 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_34_663 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.i_regbuf\[8\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[8\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[12\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_58_clk VGND VPWR clknet_3_0__leaf_clk clknet_leaf_58_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_5690_ VGND VPWR VGND VPWR _2348_ _2336_ _2341_ i_debug_uart_tx.data_to_send\[3\]
+ _2347_ sky130_fd_sc_hd__a211o_1
X_4710_ VPWR VGND _1546_ _1516_ VPWR VGND sky130_fd_sc_hd__buf_6
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.i_regbuf\[6\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[6\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[10\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_16_118 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_4641_ VPWR VGND VPWR VGND _1477_ _1473_ _1476_ sky130_fd_sc_hd__or2_2
XFILLER_0_44_449 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_71_246 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4572_ VGND VPWR VPWR VGND _1408_ _0653_ _1208_ _1407_ sky130_fd_sc_hd__mux2_4
X_7360_ VPWR VGND VGND VPWR net127 _3620_ _3619_ sky130_fd_sc_hd__nand2_1
X_6311_ VGND VPWR VPWR VGND _2766_ _2322_ _2762_ net245 sky130_fd_sc_hd__mux2_1
XFILLER_0_52_493 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_7291_ VGND VPWR _3566_ _3556_ _3555_ _3565_ VPWR VGND sky130_fd_sc_hd__and3_1
X_6242_ VPWR VGND VGND VPWR _2721_ _2719_ _2720_ sky130_fd_sc_hd__or2_1
X_6173_ VGND VPWR _1386_ _2667_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_5124_ VPWR VGND VGND VPWR _1879_ _1882_ _1881_ sky130_fd_sc_hd__nand2_1
X_5055_ VGND VPWR VPWR VGND _1812_ _1816_ _1815_ sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_49_clk VGND VPWR clknet_3_4__leaf_clk clknet_leaf_49_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_4006_ VPWR VGND VGND VPWR i_tinyqv.cpu.debug_instr_valid _0857_ i_tinyqv.cpu.is_lui
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5957_ VGND VPWR VPWR VGND _2537_ _2536_ _2524_ i_tinyqv.cpu.data_addr\[16\] sky130_fd_sc_hd__mux2_1
X_4908_ VGND VPWR VPWR VGND _1699_ _1380_ _1696_ i_tinyqv.cpu.i_core.i_registers.reg_access\[2\]\[2\]
+ sky130_fd_sc_hd__mux2_1
X_5888_ VGND VPWR _0231_ _2489_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7627_ i_tinyqv.cpu.i_core.i_registers.reg_access\[12\]\[2\] clknet_leaf_44_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[6\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.i_regbuf\[12\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[12\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[16\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4839_ VGND VPWR VPWR VGND _1660_ i_tinyqv.cpu.debug_rd\[0\] _1659_ i_tinyqv.cpu.i_core.i_registers.reg_access\[11\]\[0\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_641 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_28_490 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_7558_ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[1\] clknet_leaf_55_clk _0051_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6509_ VPWR VGND VGND VPWR _2791_ _2800_ _2918_ _2923_ sky130_fd_sc_hd__o21a_1
X_7489_ VPWR VGND VPWR VGND _3727_ _3726_ _3017_ _3728_ sky130_fd_sc_hd__a21oi_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.i_regbuf\[5\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[5\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[9\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 net93 i_tinyqv.mem.q_ctrl.addr\[1\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 net115 i_tinyqv.cpu.data_out\[22\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 net126 i_tinyqv.mem.q_ctrl.addr\[2\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 net104 i_tinyqv.cpu.i_core.i_registers.reg_access\[15\]\[2\] VPWR VGND VGND
+ VPWR sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_6 _2507_ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xrebuffer18 VGND VPWR net47 _0643_ VPWR VGND sky130_fd_sc_hd__buf_1
Xrebuffer29 VGND VPWR net58 _0645_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6860_ VGND VPWR VPWR VGND _3230_ _3229_ _3047_ _3223_ sky130_fd_sc_hd__mux2_1
X_6791_ VPWR VGND VGND VPWR i_tinyqv.cpu.instr_data_start\[16\] _3167_ i_tinyqv.cpu.imm\[16\]
+ sky130_fd_sc_hd__nand2_1
X_5811_ VPWR VGND VPWR VGND _2439_ _2437_ _2436_ _2440_ sky130_fd_sc_hd__a21oi_1
X_5742_ VGND VPWR i_spi.busy _2386_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_8530_ i_tinyqv.cpu.i_core.i_instrret.cy clknet_leaf_50_clk _0600_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_438 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_5673_ VPWR VGND VGND VPWR i_debug_uart_tx.fsm_state\[2\] i_debug_uart_tx.fsm_state\[1\]
+ i_debug_uart_tx.fsm_state\[3\] _2334_ sky130_fd_sc_hd__o21a_1
X_8461_ i_tinyqv.cpu.i_core.i_registers.rs1\[0\] clknet_leaf_51_clk _0559_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_8392_ i_tinyqv.cpu.data_out\[17\] clknet_leaf_26_clk _0490_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_7412_ VPWR VGND VGND VPWR _3662_ _3661_ _3010_ _3663_ sky130_fd_sc_hd__nor3_1
X_4624_ VGND VPWR VGND VPWR _1460_ _1408_ _1457_ _1458_ _1459_ sky130_fd_sc_hd__a22o_4
XPHY_EDGE_ROW_6_Right_6 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7343_ VPWR VGND VGND VPWR _2140_ _3607_ _3282_ _3606_ _3563_ sky130_fd_sc_hd__o211ai_1
X_4555_ VPWR VGND _1391_ _0835_ _0826_ _1388_ _1390_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_4486_ VPWR VGND VPWR VGND _0819_ _0783_ _1173_ _1325_ sky130_fd_sc_hd__a21oi_1
X_7274_ VPWR VGND VPWR VGND _3362_ _3551_ _2131_ _3552_ sky130_fd_sc_hd__or3_1
X_6225_ VPWR VGND VGND VPWR _2705_ _2702_ _2703_ sky130_fd_sc_hd__or2_1
X_6156_ VGND VPWR _0330_ _2658_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5107_ VGND VPWR VPWR VGND _1864_ _1866_ _1865_ sky130_fd_sc_hd__xor2_1
X_6087_ VGND VPWR _0308_ _2611_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5038_ VGND VPWR VPWR VGND _1797_ _1800_ _1799_ sky130_fd_sc_hd__xor2_1
X_6989_ VPWR VGND _3311_ _3310_ _3303_ _3281_ _2066_ VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_48_541 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_16_471 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_31_496 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.i_regbuf\[12\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[12\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[16\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_608 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_59_Right_59 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_10_603 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_10_625 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4340_ _1186_ _0878_ _0857_ _0858_ _1185_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
X_4271_ VPWR VGND VPWR VGND _1109_ _1092_ _1117_ _1118_ sky130_fd_sc_hd__a21oi_1
X_6010_ VGND VPWR VPWR VGND _2571_ i_tinyqv.cpu.instr_data\[2\]\[9\] _2563_ _2318_
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_68_Right_68 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7961_ i_tinyqv.cpu.i_core.mepc\[21\] clknet_leaf_35_clk _0098_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_6912_ VPWR VGND VGND VPWR _3260_ _3267_ _0772_ sky130_fd_sc_hd__nor2_2
X_7892_ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[15\] clknet_leaf_48_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[15\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6843_ VGND VPWR VGND VPWR _0461_ i_tinyqv.cpu.instr_data_start\[20\] _3123_ _3214_
+ _3205_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_77_Right_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6774_ VPWR VGND VPWR VGND i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[22\] _3039_
+ _3152_ _3151_ _3051_ _3028_ sky130_fd_sc_hd__a221o_1
X_3986_ VPWR VGND VGND VPWR i_tinyqv.cpu.no_write_in_progress _0836_ i_tinyqv.cpu.debug_instr_valid
+ _0837_ sky130_fd_sc_hd__o21a_1
XFILLER_0_45_500 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5725_ VGND VPWR VPWR VGND _2371_ i_debug_uart_tx.fsm_state\[1\] _2368_ _2372_ sky130_fd_sc_hd__or3b_1
X_8513_ i_tinyqv.cpu.i_core.i_instrret.register\[19\] clknet_leaf_45_clk i_tinyqv.cpu.i_core.i_instrret.reg_buf\[19\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5656_ VGND VPWR i_tinyqv.cpu.instr_data_in\[11\] _2322_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_8444_ i_tinyqv.cpu.imm\[22\] clknet_leaf_22_clk _0542_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4607_ VGND VPWR _0841_ _1442_ _1443_ _0653_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_5587_ VPWR VGND VGND VPWR _2272_ i_uart_rx.recieved_data\[7\] _2264_ sky130_fd_sc_hd__or2_1
X_8375_ i_debug_uart_tx.uart_tx_data\[0\] clknet_leaf_25_clk _0473_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
X_4538_ VPWR VGND VPWR VGND _1362_ _0956_ _1376_ _1377_ sky130_fd_sc_hd__a21oi_1
X_7326_ VGND VPWR _0564_ _3594_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4469_ VPWR VGND VPWR VGND _1308_ _1244_ sky130_fd_sc_hd__inv_2
X_7257_ VGND VPWR VPWR VGND _3538_ _3537_ _3395_ net69 sky130_fd_sc_hd__mux2_1
X_6208_ VGND VPWR VPWR VGND _2690_ _2688_ _2689_ debug_register_data sky130_fd_sc_hd__mux2_1
X_7188_ VGND VPWR _3486_ _3484_ _3359_ _3485_ VPWR VGND sky130_fd_sc_hd__and3_1
X_6139_ VGND VPWR _0325_ _2646_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xrebuffer9 VPWR VGND VPWR VGND net38 i_tinyqv.cpu.i_core.i_registers.rs2\[0\] sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_48_39 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_3840_ VPWR VGND VPWR VGND _0619_ i_tinyqv.cpu.imm\[15\] _0617_ _0692_ i_tinyqv.cpu.i_core.imm_lo\[7\]
+ sky130_fd_sc_hd__a22o_1
X_3771_ VPWR VGND VPWR VGND i_tinyqv.cpu.instr_data_start\[23\] _0610_ _0623_ _0613_
+ i_tinyqv.cpu.instr_data_start\[19\] _0622_ sky130_fd_sc_hd__a221o_1
X_5510_ VGND VPWR _2215_ _2200_ _2219_ i_uart_tx.cycle_counter\[9\] VPWR VGND sky130_fd_sc_hd__o21ai_1
X_6490_ VGND VPWR VPWR VGND _2905_ net274 _2897_ i_tinyqv.mem.q_ctrl.spi_in_buffer\[3\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_599 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5441_ VGND VPWR VPWR VGND _2153_ _2167_ _2164_ _2168_ sky130_fd_sc_hd__or3b_1
XFILLER_0_1_121 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5372_ VGND VPWR _2105_ i_tinyqv.cpu.i_core.imm_lo\[9\] i_tinyqv.cpu.i_core.imm_lo\[8\]
+ _1392_ VPWR VGND sky130_fd_sc_hd__and3_1
X_8160_ i_tinyqv.cpu.instr_data\[2\]\[9\] clknet_leaf_10_clk _0272_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_8091_ gpio_out\[2\] clknet_leaf_19_clk _0002_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4323_ VPWR VGND VPWR VGND _1170_ _0847_ sky130_fd_sc_hd__inv_2
X_7111_ VPWR VGND VPWR VGND _3363_ _2165_ _3351_ _3419_ _3418_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_198 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_7042_ VPWR VGND VGND VPWR _1468_ _3306_ _1456_ _3355_ _3356_ sky130_fd_sc_hd__o22a_1
X_4254_ VGND VPWR VPWR VGND _1101_ i_tinyqv.cpu.i_core.i_shift.a\[8\] _1028_ i_tinyqv.cpu.i_core.i_shift.a\[23\]
+ sky130_fd_sc_hd__mux2_1
X_4185_ VPWR VGND VPWR VGND _0844_ _1031_ i_tinyqv.cpu.alu_op\[3\] _1030_ _1032_ sky130_fd_sc_hd__or4_1
X_7944_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[3\] clknet_leaf_50_clk _0057_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7875_ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[30\] clknet_leaf_3_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[30\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6826_ VGND VPWR VPWR VGND _3197_ _3199_ _3198_ sky130_fd_sc_hd__xor2_1
X_6757_ VPWR VGND VGND VPWR i_tinyqv.cpu.instr_data_start\[13\] _3136_ i_tinyqv.cpu.imm\[13\]
+ sky130_fd_sc_hd__nand2_1
X_5708_ VPWR VGND VPWR VGND _2356_ _2358_ _2359_ _0182_ sky130_fd_sc_hd__a21oi_1
X_3969_ VGND VPWR VGND VPWR _0821_ _0820_ _0819_ _0783_ _0817_ sky130_fd_sc_hd__o211ai_2
X_6688_ VGND VPWR VPWR VGND _3073_ _3072_ _2987_ _1593_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_599 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_8427_ i_tinyqv.cpu.i_core.imm_lo\[5\] clknet_leaf_9_clk _0525_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_5_460 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.i_regbuf\[30\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[30\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[2\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5639_ VGND VPWR VPWR VGND _2312_ i_tinyqv.cpu.instr_data_in\[4\] _2309_ i_tinyqv.cpu.instr_data\[3\]\[4\]
+ sky130_fd_sc_hd__mux2_1
X_8358_ i_tinyqv.cpu.instr_data_start\[16\] clknet_leaf_36_clk _0457_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
X_7309_ VPWR VGND VPWR VGND _1468_ _3580_ _3581_ _3572_ _1501_ _3497_ sky130_fd_sc_hd__a221o_1
Xhold150 net179 i_tinyqv.cpu.i_core.mie\[18\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_591 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold161 net190 i_tinyqv.cpu.imm\[26\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 net201 i_uart_rx.recieved_data\[1\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_8289_ i_tinyqv.mem.qspi_data_buf\[29\] clknet_leaf_14_clk _0388_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
Xhold183 net212 i_tinyqv.cpu.is_lui VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 net223 i_tinyqv.cpu.i_core.mepc\[22\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.i_regbuf\[26\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[26\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[30\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_19 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.i_regbuf\[15\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[15\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[19\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_580 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_75_37 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_instrret.i_regbuf\[25\] i_tinyqv.cpu.i_core.i_instrret.reg_buf\[25\]
+ i_tinyqv.cpu.i_core.i_instrret.register\[29\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5990_ VPWR VGND VPWR VGND _2552_ i_tinyqv.cpu.data_addr\[27\] _1758_ _2559_ i_tinyqv.cpu.i_core.i_shift.a\[31\]
+ sky130_fd_sc_hd__a22o_1
X_4941_ VPWR VGND VGND VPWR _1723_ _1716_ _1722_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_425 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4872_ VGND VPWR VPWR VGND _1678_ net32 _1674_ i_tinyqv.cpu.i_core.i_registers.reg_access\[8\]\[3\]
+ sky130_fd_sc_hd__mux2_1
X_7660_ i_tinyqv.cpu.i_core.i_registers.reg_access\[11\]\[3\] clknet_leaf_45_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[7\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6611_ VGND VPWR _3006_ _3007_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_3823_ VGND VPWR VGND VPWR _0663_ _0675_ i_tinyqv.cpu.i_core.i_registers.rs2\[2\]
+ net38 i_tinyqv.cpu.i_core.i_registers.rs2\[3\] sky130_fd_sc_hd__and4bb_2
X_7591_ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[2\] clknet_leaf_55_clk _0048_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6542_ VPWR VGND _2952_ _2916_ _1713_ VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_15_536 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_27_396 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_6473_ VGND VPWR VPWR VGND _0410_ _2895_ _2894_ _2629_ _2596_ i_tinyqv.cpu.i_core.i_shift.a\[29\]
+ sky130_fd_sc_hd__a32o_1
X_8212_ i_tinyqv.cpu.instr_data\[0\]\[1\] clknet_leaf_13_clk _0324_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5424_ VGND VPWR VPWR VGND _2154_ i_tinyqv.cpu.i_core.i_registers.rd\[0\] _2153_
+ _2148_ sky130_fd_sc_hd__mux2_1
X_8143_ i_tinyqv.cpu.data_addr\[18\] clknet_leaf_34_clk _0255_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_452 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_57_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5355_ VPWR VGND VPWR VGND _2090_ _0729_ _2056_ _2092_ _2091_ sky130_fd_sc_hd__a22o_1
X_5286_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[14\] _2038_ _1845_ sky130_fd_sc_hd__nand2_1
X_4306_ VGND VPWR VGND VPWR _1153_ _1120_ _1091_ _1149_ _1152_ sky130_fd_sc_hd__a211o_1
X_8074_ i_tinyqv.cpu.i_core.mie\[17\] clknet_leaf_37_clk _0209_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_4237_ VGND VPWR VPWR VGND _1084_ _1082_ _1083_ _1081_ sky130_fd_sc_hd__mux2_1
X_7025_ VPWR VGND VGND VPWR _1490_ _1494_ _3341_ sky130_fd_sc_hd__nor2_1
X_4168_ VPWR VGND VPWR VGND _1015_ _0866_ sky130_fd_sc_hd__inv_2
X_4099_ VPWR VGND VGND VPWR _0946_ _0908_ _0945_ sky130_fd_sc_hd__nand2_2
X_7927_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[18\] clknet_leaf_25_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[18\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7858_ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[13\] clknet_leaf_47_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[13\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6809_ VPWR VGND VGND VPWR _3037_ _3184_ _3183_ sky130_fd_sc_hd__nand2_1
X_7789_ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[8\] clknet_leaf_2_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[8\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.i_regbuf\[31\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[31\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[3\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_672 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.i_regbuf\[27\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[27\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[31\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.i_regbuf\[16\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[16\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[20\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_296 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.i_regbuf\[30\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[30\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[2\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_697 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5140_ VPWR VGND VGND VPWR _1898_ _1894_ _1896_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_594 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_5071_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[5\] _1831_ _1789_ sky130_fd_sc_hd__nand2_1
X_4022_ VPWR VGND VGND VPWR _0871_ _0870_ _0867_ _0872_ sky130_fd_sc_hd__nor3_1
X_5973_ VGND VPWR _0258_ _2547_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4924_ VPWR VGND VGND VPWR _1709_ _1708_ _1706_ sky130_fd_sc_hd__nor2_4
X_7712_ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[27\] clknet_leaf_59_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[27\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4855_ VGND VPWR _0033_ _1668_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7643_ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[22\] clknet_leaf_46_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[22\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4786_ VGND VPWR VPWR VGND _1621_ i_tinyqv.mem.qspi_data_buf\[15\] _1017_ i_tinyqv.cpu.instr_data_in\[15\]
+ sky130_fd_sc_hd__mux2_1
X_7574_ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[17\] clknet_leaf_58_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[17\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_3806_ VGND VPWR _0657_ _0658_ VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_6525_ VGND VPWR VPWR VGND _2937_ i_tinyqv.cpu.data_out\[18\] _2911_ i_tinyqv.cpu.data_out\[26\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_491 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_15_388 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_43_664 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_6456_ VPWR VGND _2882_ _2855_ _2810_ i_tinyqv.mem.q_ctrl.spi_clk_out _2881_ VGND
+ VPWR sky130_fd_sc_hd__a31o_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.i_regbuf\[9\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[9\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[13\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6387_ VPWR VGND _2826_ _2783_ _2790_ i_tinyqv.mem.q_ctrl.delay_cycles_cfg\[2\] _2825_
+ VGND VPWR sky130_fd_sc_hd__a31o_1
X_5407_ VPWR VGND VPWR VGND _2134_ _2136_ _2121_ _2137_ sky130_fd_sc_hd__or3_1
X_8126_ i_tinyqv.cpu.data_addr\[1\] clknet_leaf_33_clk _0238_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5338_ VPWR VGND VGND VPWR _2077_ _2078_ _0093_ sky130_fd_sc_hd__nor2_1
X_8057_ i_spi.data\[0\] clknet_leaf_27_clk _0192_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5269_ VGND VPWR VPWR VGND _2019_ _0017_ _2021_ sky130_fd_sc_hd__xor2_1
X_7008_ VGND VPWR VPWR VGND _3327_ _3326_ _3281_ i_tinyqv.cpu.is_alu_reg sky130_fd_sc_hd__mux2_1
XFILLER_0_65_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_18_160 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_25_108 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_1_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_33_174 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_16 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.i_regbuf\[8\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[8\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[12\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_4640_ VGND VPWR VPWR VGND _1476_ _1408_ _1475_ _1474_ sky130_fd_sc_hd__mux2_4
X_6310_ VGND VPWR _0377_ _2765_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4571_ VPWR VGND VPWR VGND _1407_ _0749_ sky130_fd_sc_hd__inv_2
X_7290_ VPWR VGND VPWR VGND _2165_ _3305_ _3287_ _3565_ sky130_fd_sc_hd__a21oi_1
X_6241_ VGND VPWR _2720_ _2715_ _2698_ _2718_ VPWR VGND sky130_fd_sc_hd__and3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.i_regbuf\[20\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[20\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[24\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6172_ VGND VPWR _0338_ _2666_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.i_regbuf\[6\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[6\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[10\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5123_ VPWR VGND VPWR VGND _1789_ _1054_ _1880_ _1881_ i_tinyqv.cpu.i_core.i_shift.a\[6\]
+ sky130_fd_sc_hd__a22o_1
X_5054_ VPWR VGND _1815_ _1813_ _1767_ i_tinyqv.cpu.i_core.i_shift.a\[3\] _1814_ VGND
+ VPWR sky130_fd_sc_hd__a31o_1
X_4005_ _0856_ _0854_ _0852_ _0853_ _0855_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
XFILLER_0_48_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_5956_ VGND VPWR VPWR VGND _2536_ i_tinyqv.cpu.i_core.mepc\[16\] _2504_ i_tinyqv.cpu.i_core.i_shift.a\[20\]
+ sky130_fd_sc_hd__mux2_1
X_5887_ VGND VPWR VPWR VGND _2489_ _2488_ _2399_ i_spi.data\[2\] sky130_fd_sc_hd__mux2_1
X_4907_ VGND VPWR _0059_ _1698_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7626_ i_tinyqv.cpu.i_core.i_registers.reg_access\[12\]\[1\] clknet_leaf_55_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[5\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4838_ i_tinyqv.cpu.i_core.i_registers.rd\[0\] _1659_ i_tinyqv.cpu.i_core.i_registers.rd\[1\]
+ _1658_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_7557_ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[0\] clknet_leaf_53_clk _0050_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_686 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_4769_ VGND VPWR _0841_ _1604_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_6508_ VGND VPWR VPWR VGND _2922_ _2921_ _2792_ _2917_ sky130_fd_sc_hd__mux2_1
X_7488_ VPWR VGND VGND VPWR _3727_ i_tinyqv.cpu.instr_data_start\[22\] _3720_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_494 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6439_ VPWR VGND VPWR VGND _2869_ _2870_ _2853_ _2871_ _2863_ sky130_fd_sc_hd__or4b_1
XFILLER_0_30_188 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_8109_ i_tinyqv.cpu.instr_data\[0\]\[9\] clknet_leaf_10_clk _0221_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
Xhold65 net94 i_tinyqv.cpu.data_continue VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 net116 i_uart_tx.data_to_send\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 net127 i_tinyqv.cpu.i_core.is_interrupt VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 net105 i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[24\] VPWR VGND VGND
+ VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.i_regbuf\[5\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[5\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[9\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_704 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_53_236 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_38_299 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XANTENNA_7 _2734_ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_0_22_645 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xrebuffer19 VGND VPWR net48 net47 VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5810_ VGND VPWR VGND VPWR _2439_ _2438_ _0613_ i_tinyqv.cpu.i_core.interrupt_req\[1\]
+ i_tinyqv.cpu.i_core.mip\[17\] sky130_fd_sc_hd__a211o_1
X_6790_ VPWR VGND VGND VPWR _3166_ i_tinyqv.cpu.instr_data_start\[16\] i_tinyqv.cpu.imm\[16\]
+ sky130_fd_sc_hd__or2_1
XFILLER_0_9_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_5741_ VPWR VGND VGND VPWR i_spi.busy _2385_ i_spi.clock_count\[0\] sky130_fd_sc_hd__nand2_1
XFILLER_0_8_149 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_8460_ i_tinyqv.cpu.i_core.mem_op\[2\] clknet_leaf_7_clk _0558_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_5672_ VPWR VGND _2333_ _2332_ VPWR VGND sky130_fd_sc_hd__buf_2
X_7411_ VPWR VGND VPWR VGND _3651_ _0882_ i_tinyqv.cpu.instr_data_start\[10\] _3662_
+ sky130_fd_sc_hd__a21oi_1
X_8391_ i_tinyqv.cpu.data_out\[16\] clknet_leaf_26_clk _0489_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_4623_ VGND VPWR VPWR VGND _1459_ i_tinyqv.cpu.instr_data\[2\]\[2\] _1412_ i_tinyqv.cpu.instr_data\[0\]\[2\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_645 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7342_ VPWR VGND VPWR VGND _1510_ _2143_ _3606_ _3351_ _1460_ _3328_ sky130_fd_sc_hd__a221o_1
X_4554_ VPWR VGND VGND VPWR i_tinyqv.cpu.is_branch _1390_ _0653_ sky130_fd_sc_hd__nand2_4
X_7273_ VGND VPWR VPWR VGND _3551_ _3549_ _3531_ _3467_ _3550_ _2121_ sky130_fd_sc_hd__a32o_1
X_6224_ VPWR VGND VGND VPWR _2702_ _2704_ _2703_ sky130_fd_sc_hd__nand2_1
X_4485_ VPWR VGND VGND VPWR _1324_ _0783_ _0819_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_6155_ VGND VPWR VPWR VGND _2658_ net264 _2656_ i_tinyqv.cpu.i_core.mepc\[1\] sky130_fd_sc_hd__mux2_1
X_5106_ VGND VPWR VGND VPWR _1865_ _1840_ i_tinyqv.cpu.i_core.multiplier.accum\[7\]
+ _1838_ sky130_fd_sc_hd__a21bo_1
X_6086_ VGND VPWR VPWR VGND _2611_ _1060_ _2596_ i_tinyqv.cpu.i_core.i_shift.a\[19\]
+ sky130_fd_sc_hd__mux2_1
X_5037_ VPWR VGND VPWR VGND _1774_ i_tinyqv.cpu.i_core.multiplier.accum\[4\] _1798_
+ _1799_ sky130_fd_sc_hd__a21o_1
X_6988_ _3310_ _3304_ _3305_ _3306_ _3309_ VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_5939_ VGND VPWR VPWR VGND _2525_ _2523_ _2524_ i_tinyqv.cpu.data_addr\[10\] sky130_fd_sc_hd__mux2_1
XFILLER_0_35_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_7609_ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[20\] clknet_leaf_0_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[20\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.i_regbuf\[20\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[20\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[24\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_589 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4270_ VPWR VGND VPWR VGND _1116_ _1080_ _1076_ _1117_ sky130_fd_sc_hd__a21o_1
X_7960_ i_tinyqv.cpu.i_core.mepc\[20\] clknet_leaf_36_clk _0097_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_6911_ VGND VPWR VPWR VGND _0477_ _3265_ _3261_ _1619_ _3266_ net309 sky130_fd_sc_hd__a32o_1
X_7891_ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[14\] clknet_leaf_2_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[14\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6842_ VPWR VGND VGND VPWR _3214_ _3029_ _3213_ sky130_fd_sc_hd__or2_1
X_6773_ VGND VPWR VPWR VGND _3151_ _3150_ _2991_ _2532_ sky130_fd_sc_hd__mux2_1
X_3985_ VPWR VGND VGND VPWR i_tinyqv.cpu.is_store i_tinyqv.cpu.is_load _0836_ sky130_fd_sc_hd__nor2_1
X_5724_ VPWR VGND VGND VPWR _2339_ _2333_ _2371_ sky130_fd_sc_hd__nor2_1
X_8512_ i_tinyqv.cpu.i_core.i_instrret.register\[18\] clknet_leaf_49_clk i_tinyqv.cpu.i_core.i_instrret.reg_buf\[18\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5655_ VGND VPWR _0167_ _2321_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8443_ i_tinyqv.cpu.imm\[21\] clknet_leaf_7_clk _0541_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_8374_ i_tinyqv.cpu.load_started clknet_leaf_21_clk _0472_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4606_ VPWR VGND _1442_ _1441_ VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_0_4_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5586_ VGND VPWR VGND VPWR _0148_ net172 _2263_ _2271_ _2240_ sky130_fd_sc_hd__o211a_1
XFILLER_0_13_442 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_7325_ VGND VPWR VPWR VGND _3594_ _0663_ _2153_ _3593_ sky130_fd_sc_hd__mux2_1
X_4537_ VPWR VGND VGND VPWR _0957_ _1369_ _0982_ _1375_ _1376_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_15_Left_96 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_40_272 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_4468_ VGND VPWR _1307_ uo_out[6] VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_7256_ VGND VPWR VGND VPWR _3537_ _3534_ _3536_ _3531_ _2129_ sky130_fd_sc_hd__a211o_1
X_6207_ VPWR VGND _2689_ _0995_ _0970_ _0984_ _2198_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_7187_ VGND VPWR VGND VPWR _3485_ _3331_ _3471_ _3304_ _3481_ sky130_fd_sc_hd__a211o_1
X_4399_ VPWR VGND VPWR VGND _1223_ _0956_ _1241_ _1242_ sky130_fd_sc_hd__a21o_1
X_6138_ VGND VPWR VPWR VGND _2646_ _2644_ _2645_ _1083_ sky130_fd_sc_hd__mux2_1
X_6069_ VGND VPWR _0299_ _2602_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_3770_ VPWR VGND VGND VPWR _0618_ _0621_ _0611_ _0622_ sky130_fd_sc_hd__o21a_1
X_5440_ VPWR VGND VPWR VGND _2121_ _2166_ _2141_ _2149_ _2167_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_5371_ VGND VPWR VPWR VGND _2104_ _2103_ _2057_ i_tinyqv.cpu.i_core.mstatus_mie sky130_fd_sc_hd__mux2_1
X_8090_ gpio_out\[1\] clknet_leaf_27_clk _0001_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4322_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[0\] i_tinyqv.cpu.i_core.multiplier.accum\[0\]
+ _1169_ _1167_ sky130_fd_sc_hd__nand3_1
X_7110_ VPWR VGND VGND VPWR _3368_ i_tinyqv.cpu.instr_data\[1\]\[9\] _3366_ i_tinyqv.cpu.instr_data\[0\]\[9\]
+ _3418_ _3417_ sky130_fd_sc_hd__o221a_1
XFILLER_0_1_177 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4253_ VPWR VGND VGND VPWR _1092_ _1100_ _1099_ sky130_fd_sc_hd__nand2_1
X_7041_ VPWR VGND VGND VPWR _3355_ _3348_ _3354_ sky130_fd_sc_hd__or2_1
X_4184_ VGND VPWR VGND VPWR _0842_ i_tinyqv.cpu.i_core.cycle\[1\] _1031_ sky130_fd_sc_hd__or2_4
X_7943_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[2\] clknet_leaf_50_clk _0056_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7874_ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[29\] clknet_leaf_47_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[29\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6825_ VGND VPWR _3186_ _3188_ _3198_ _3187_ VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_211 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6756_ VGND VPWR _2987_ _3134_ _3135_ _1201_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_3968_ VPWR VGND VGND VPWR net80 _0820_ _0700_ sky130_fd_sc_hd__nand2_1
X_5707_ VGND VPWR _2356_ _2357_ _2359_ _2358_ VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_578 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_3899_ VPWR VGND VPWR VGND i_tinyqv.cpu.instr_data_start\[5\] _0748_ _0751_ _0690_
+ i_tinyqv.cpu.instr_data_start\[9\] _0750_ sky130_fd_sc_hd__a221o_1
X_6687_ VPWR VGND VPWR VGND _3072_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[15\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_60_334 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5638_ VGND VPWR _0160_ _2311_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8426_ i_tinyqv.cpu.i_core.imm_lo\[4\] clknet_leaf_9_clk _0524_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_2
X_5569_ VPWR VGND VPWR VGND _2259_ net142 _2261_ _0141_ sky130_fd_sc_hd__a21oi_1
X_8357_ i_tinyqv.cpu.instr_data_start\[15\] clknet_leaf_36_clk _0456_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.i_regbuf\[23\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[23\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[27\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 net191 i_uart_rx.bit_sample VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold140 net169 i_spi.dc_in VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 net180 i_tinyqv.cpu.data_ready_latch VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7308_ VPWR VGND VGND VPWR _1473_ _3321_ _3580_ sky130_fd_sc_hd__nor2_1
Xhold195 net224 i_uart_rx.cycle_counter\[2\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 net202 _0142_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_8288_ i_tinyqv.mem.qspi_data_buf\[28\] clknet_leaf_14_clk _0387_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
Xhold184 net213 i_tinyqv.cpu.imm\[16\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7239_ VPWR VGND _3524_ _3441_ _3330_ _3291_ _3510_ VGND VPWR sky130_fd_sc_hd__a31o_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.i_regbuf\[19\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[19\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[23\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_209 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xi_tinyqv.cpu.i_core.i_instrret.i_regbuf\[18\] i_tinyqv.cpu.i_core.i_instrret.reg_buf\[18\]
+ i_tinyqv.cpu.i_core.i_instrret.register\[22\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4940_ VPWR VGND VPWR VGND _1706_ _1721_ _1722_ i_tinyqv.mem.q_ctrl.addr\[23\] _1709_
+ _1719_ sky130_fd_sc_hd__a221o_1
X_4871_ VGND VPWR _0076_ _1677_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6610_ VPWR VGND i_tinyqv.mem.q_ctrl.spi_clk_out _3006_ _1709_ VPWR VGND sky130_fd_sc_hd__and2_2
X_7590_ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[1\] clknet_leaf_55_clk _0047_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_3822_ VGND VPWR VGND VPWR net38 _0674_ i_tinyqv.cpu.i_core.i_registers.rs2\[2\]
+ i_tinyqv.cpu.i_core.i_registers.rs2\[3\] net37 sky130_fd_sc_hd__and4bb_2
X_6541_ VGND VPWR _0422_ _2951_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_651 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6472_ VPWR VGND VGND VPWR net66 _2895_ _0845_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_323 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_8211_ i_tinyqv.cpu.instr_data\[0\]\[0\] clknet_leaf_9_clk _0323_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5423_ VPWR VGND VGND VPWR _2152_ _2153_ _1752_ sky130_fd_sc_hd__nand2_4
X_8142_ i_tinyqv.cpu.data_addr\[17\] clknet_leaf_34_clk _0254_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_5354_ VPWR VGND VPWR VGND net18 _1312_ _2056_ _2091_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4305_ VPWR VGND VGND VPWR _1088_ _1151_ _1152_ sky130_fd_sc_hd__nor2_1
X_5285_ VPWR VGND VGND VPWR _2035_ _2037_ _2036_ sky130_fd_sc_hd__nand2_1
X_8073_ i_tinyqv.cpu.i_core.mie\[18\] clknet_leaf_38_clk _0208_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_4236_ VGND VPWR _1050_ _1083_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_7024_ VPWR VGND _3340_ _3295_ i_tinyqv.cpu.is_jalr VPWR VGND sky130_fd_sc_hd__and2_1
X_4167_ VGND VPWR VPWR VGND _1014_ i_tinyqv.mem.qspi_data_buf\[12\] _0838_ i_tinyqv.mem.qspi_data_buf\[8\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_27_Left_108 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4098_ VPWR VGND VGND VPWR _0907_ _0945_ _0688_ sky130_fd_sc_hd__nor2_2
X_7926_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[17\] clknet_leaf_25_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[17\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7857_ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[12\] clknet_leaf_49_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[12\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6808_ VPWR VGND VPWR VGND _3174_ _3039_ _3183_ _2306_ _1213_ _3182_ sky130_fd_sc_hd__a221o_1
X_7788_ i_tinyqv.cpu.i_core.i_registers.reg_access\[7\]\[3\] clknet_leaf_1_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[7\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6739_ VGND VPWR VPWR VGND _3120_ _3119_ _2990_ _2526_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_36_Left_117 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.i_regbuf\[24\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[24\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[28\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_8409_ VGND VPWR VGND VPWR i_tinyqv.cpu.counter\[4\] _0507_ clknet_leaf_22_clk sky130_fd_sc_hd__dfxtp_4
XPHY_EDGE_ROW_45_Left_126 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_29_629 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_54_Left_135 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_37_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.i_regbuf\[23\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[23\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[27\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_518 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_cycles.i_regbuf\[21\] i_tinyqv.cpu.i_core.i_cycles.reg_buf\[21\]
+ i_tinyqv.cpu.i_core.i_cycles.register\[25\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_63_Left_144 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.i_regbuf\[12\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[12\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[16\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5070_ _1830_ _1824_ _1822_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_4021_ VPWR VGND VGND VPWR _0868_ _0869_ _0871_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_52 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5972_ VGND VPWR VPWR VGND _2547_ _2546_ _2501_ i_tinyqv.cpu.data_addr\[21\] sky130_fd_sc_hd__mux2_1
X_4923_ VPWR VGND VGND VPWR _1707_ i_tinyqv.mem.q_ctrl.fsm_state\[1\] _1708_ sky130_fd_sc_hd__or2b_2
X_7711_ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[26\] clknet_leaf_52_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[26\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_72_Left_153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_51_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4854_ VGND VPWR VPWR VGND _1668_ i_tinyqv.cpu.debug_rd\[3\] _1664_ i_tinyqv.cpu.i_core.i_registers.reg_access\[10\]\[3\]
+ sky130_fd_sc_hd__mux2_1
X_7642_ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[21\] clknet_leaf_55_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[21\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4785_ VGND VPWR VGND VPWR _1620_ _0957_ _1615_ _1618_ _1619_ sky130_fd_sc_hd__o211a_1
X_7573_ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[16\] clknet_leaf_59_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[16\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_556 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_7_545 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_3805_ VPWR VGND VGND VPWR _0657_ _0656_ i_tinyqv.cpu.alu_op\[3\] sky130_fd_sc_hd__or2_1
X_6524_ VGND VPWR VPWR VGND _2936_ i_tinyqv.cpu.data_out\[10\] _2909_ i_debug_uart_tx.uart_tx_data\[2\]
+ sky130_fd_sc_hd__mux2_1
X_6455_ VPWR VGND VGND VPWR i_tinyqv.mem.q_ctrl.spi_clk_out _2836_ _2881_ sky130_fd_sc_hd__nor2_1
X_6386_ VPWR VGND VPWR VGND _2825_ _2804_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_261 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_5406_ VGND VPWR _2135_ _1427_ _2136_ _1490_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_8125_ i_tinyqv.cpu.data_addr\[0\] clknet_leaf_29_clk _0237_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_5337_ VGND VPWR _2075_ _2049_ _2078_ net218 VPWR VGND sky130_fd_sc_hd__o21ai_1
X_8056_ i_spi.clock_count\[1\] clknet_leaf_27_clk _0191_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5268_ VPWR VGND VGND VPWR _1993_ _2021_ _2020_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_92 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_4219_ VGND VPWR VPWR VGND _1066_ _1065_ _1050_ _1064_ sky130_fd_sc_hd__mux2_1
X_7007_ VGND VPWR VGND VPWR _3326_ _3301_ _2136_ _2121_ _2131_ sky130_fd_sc_hd__a211o_1
X_5199_ VGND VPWR VPWR VGND _1952_ _1954_ _1953_ sky130_fd_sc_hd__xor2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.i_regbuf\[9\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[9\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[13\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7909_ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[0\] clknet_leaf_48_clk _0058_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_440 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_21_304 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_3_Left_84 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_69_584 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4570_ VPWR VGND _1406_ i_tinyqv.cpu.instr_write_offset\[1\] VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_0_52_440 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6240_ VPWR VGND VPWR VGND _2715_ _2698_ _2718_ _2719_ sky130_fd_sc_hd__a21oi_1
X_6171_ VGND VPWR VPWR VGND _2666_ net226 _2656_ i_tinyqv.cpu.i_core.mepc\[9\] sky130_fd_sc_hd__mux2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.i_regbuf\[13\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[13\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[17\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5122_ VPWR VGND _1880_ _1309_ VPWR VGND sky130_fd_sc_hd__buf_2
X_5053_ VPWR VGND VGND VPWR _1791_ _1792_ _1814_ sky130_fd_sc_hd__nor2_1
X_4004_ VPWR VGND VGND VPWR _0855_ i_tinyqv.cpu.debug_instr_valid i_tinyqv.cpu.is_system
+ sky130_fd_sc_hd__nand2_2
X_5955_ VGND VPWR _0252_ _2535_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5886_ VGND VPWR VPWR VGND _2488_ i_spi.data\[1\] _2386_ i_debug_uart_tx.uart_tx_data\[2\]
+ sky130_fd_sc_hd__mux2_1
X_4906_ VGND VPWR VPWR VGND _1698_ _1303_ _1696_ i_tinyqv.cpu.i_core.i_registers.reg_access\[2\]\[1\]
+ sky130_fd_sc_hd__mux2_1
X_7625_ i_tinyqv.cpu.i_core.i_registers.reg_access\[12\]\[0\] clknet_leaf_52_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[4\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4837_ i_tinyqv.cpu.i_core.i_registers.rd\[2\] i_tinyqv.cpu.i_core.i_registers.rd\[3\]
+ _1658_ _1188_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_7556_ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[31\] clknet_leaf_46_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[31\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_665 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_4768_ VPWR VGND VPWR VGND _1602_ _1598_ _0858_ _1603_ sky130_fd_sc_hd__a21o_1
X_6507_ VGND VPWR VPWR VGND _2921_ _2919_ _2920_ net10 sky130_fd_sc_hd__mux2_1
X_4699_ VPWR VGND VPWR VGND _1535_ _1518_ sky130_fd_sc_hd__inv_2
X_7487_ VPWR VGND VGND VPWR i_tinyqv.cpu.instr_data_start\[22\] _3726_ _3720_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_101 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_31_646 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6438_ VPWR VGND VGND VPWR i_tinyqv.mem.q_ctrl.delay_cycles_cfg\[2\] i_tinyqv.mem.q_ctrl.delay_cycles_cfg\[1\]
+ _2788_ _2870_ sky130_fd_sc_hd__o21a_1
Xi_tinyqv.cpu.i_core.i_instrret.i_regbuf\[7\] i_tinyqv.cpu.i_core.i_instrret.reg_buf\[7\]
+ i_tinyqv.cpu.i_core.i_instrret.register\[11\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_668 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6369_ VPWR VGND VPWR VGND _2810_ _1540_ sky130_fd_sc_hd__inv_2
X_8108_ i_tinyqv.cpu.instr_data\[0\]\[8\] clknet_leaf_11_clk _0220_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_370 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_8039_ i_debug_uart_tx.data_to_send\[1\] clknet_leaf_29_clk _0174_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
Xhold88 VGND VPWR i_debug_uart_tx.uart_tx_data\[0\] net117 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xhold66 net95 i_tinyqv.mem.q_ctrl.addr\[3\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 net106 i_tinyqv.cpu.instr_data\[3\]\[1\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 net128 _0029_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_8 _2930_ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_0_1_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_381 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_9_607 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_5740_ VPWR VGND VGND VPWR i_spi.busy _2384_ _2383_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_629 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_32_42 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_5671_ VGND VPWR _2332_ i_debug_uart_tx.cycle_counter\[0\] i_debug_uart_tx.cycle_counter\[2\]
+ _2331_ VPWR VGND sky130_fd_sc_hd__and3_1
X_7410_ VGND VPWR _3661_ _0882_ i_tinyqv.cpu.instr_data_start\[10\] _3651_ VPWR VGND
+ sky130_fd_sc_hd__and3_1
X_8390_ i_tinyqv.cpu.data_out\[15\] clknet_leaf_20_clk _0488_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_4622_ VPWR VGND VGND VPWR i_tinyqv.cpu.instr_data\[1\]\[2\] _1414_ _1416_ _1458_
+ sky130_fd_sc_hd__o21a_1
X_4553_ VPWR VGND VPWR VGND _0835_ _0826_ _1388_ _1389_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_7341_ VGND VPWR VGND VPWR _0568_ _3295_ _3333_ net196 _2067_ sky130_fd_sc_hd__a211o_1
X_4484_ VPWR VGND VGND VPWR _1323_ _1320_ _1321_ sky130_fd_sc_hd__or2_1
X_7272_ VGND VPWR VGND VPWR _3550_ _3288_ _2165_ _3545_ sky130_fd_sc_hd__a21bo_1
X_6223_ VPWR VGND VPWR VGND _2030_ _2028_ _2033_ _2703_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_6154_ VGND VPWR _0329_ _2657_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5105_ VPWR VGND VGND VPWR _1862_ _1864_ _1863_ sky130_fd_sc_hd__nand2_1
X_6085_ VGND VPWR _0307_ _2610_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5036_ VPWR VGND _1798_ _1773_ _1771_ VPWR VGND sky130_fd_sc_hd__and2_1
X_6987_ VPWR VGND VGND VPWR _2126_ _3309_ _3308_ sky130_fd_sc_hd__nand2_1
X_5938_ VGND VPWR _2501_ _2524_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_63_557 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5869_ VGND VPWR VPWR VGND _2479_ i_tinyqv.cpu.instr_data\[0\]\[11\] _2469_ _2322_
+ sky130_fd_sc_hd__mux2_1
X_7608_ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[19\] clknet_leaf_2_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[19\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_194 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7539_ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[14\] clknet_leaf_45_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[14\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.i_regbuf\[13\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[13\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[17\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_465 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_12_690 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_41_218 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_22_421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_6910_ VPWR VGND VGND VPWR _3266_ _0939_ _0854_ sky130_fd_sc_hd__or2_1
X_7890_ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[13\] clknet_leaf_5_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[13\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6841_ VGND VPWR VPWR VGND _3213_ _3212_ _3047_ _3206_ sky130_fd_sc_hd__mux2_1
X_6772_ VGND VPWR _3149_ _3150_ _3146_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_8511_ i_tinyqv.cpu.i_core.i_instrret.register\[17\] clknet_leaf_45_clk i_tinyqv.cpu.i_core.i_instrret.reg_buf\[17\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_3984_ VPWR VGND VGND VPWR _0826_ i_tinyqv.cpu.i_core.cmp_out _0835_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_513 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5723_ VGND VPWR VPWR VGND _0186_ _2370_ _2369_ _2221_ _2357_ i_debug_uart_tx.fsm_state\[0\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_5_610 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_259 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5654_ VGND VPWR VPWR VGND _2321_ _2320_ _2309_ i_tinyqv.cpu.instr_data\[3\]\[10\]
+ sky130_fd_sc_hd__mux2_1
X_8442_ i_tinyqv.cpu.imm\[20\] clknet_leaf_7_clk _0540_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_60_538 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_8373_ i_tinyqv.cpu.no_write_in_progress clknet_leaf_22_clk _0471_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
X_4605_ VPWR VGND VGND VPWR _1441_ _1439_ _1440_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_229 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5585_ VPWR VGND VGND VPWR _2271_ i_uart_rx.recieved_data\[6\] _2264_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_153 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7324_ VGND VPWR VPWR VGND _3593_ _3592_ _2149_ _3590_ sky130_fd_sc_hd__mux2_1
X_4536_ VPWR VGND VGND VPWR _0724_ _1370_ _1374_ _1375_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_13_465 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_13_476 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_4467_ VGND VPWR VPWR VGND _1307_ gpio_out\[6\] gpio_out_sel\[6\] i_debug_uart_tx.txd_reg
+ sky130_fd_sc_hd__mux2_1
X_7255_ VPWR VGND VPWR VGND _3535_ _3536_ _1456_ _3301_ sky130_fd_sc_hd__a21boi_1
X_6206_ VGND VPWR VPWR VGND _2688_ i_debug_uart_tx.uart_tx_data\[0\] _1728_ net5 sky130_fd_sc_hd__mux2_1
X_4398_ VPWR VGND VGND VPWR _0957_ _1234_ _0982_ _1240_ _1241_ sky130_fd_sc_hd__o22a_1
X_7186_ VPWR VGND VPWR VGND _3476_ _1486_ _3479_ _3484_ sky130_fd_sc_hd__a21o_1
X_6137_ VPWR VGND VGND VPWR _1755_ _2645_ _1026_ sky130_fd_sc_hd__nor2_2
X_6068_ VGND VPWR VPWR VGND _2602_ i_tinyqv.cpu.i_core.i_shift.a\[10\] _2593_ i_tinyqv.cpu.i_core.i_shift.a\[6\]
+ sky130_fd_sc_hd__mux2_1
X_5019_ VGND VPWR _1781_ _1578_ _1782_ _1579_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_51_505 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_64_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_39_384 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_2_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_5370_ _2103_ _2102_ net41 VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
XFILLER_0_10_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_4321_ VPWR VGND VPWR VGND _1167_ i_tinyqv.cpu.i_core.i_shift.a\[0\] i_tinyqv.cpu.i_core.multiplier.accum\[0\]
+ _1168_ sky130_fd_sc_hd__a21o_1
X_4252_ VGND VPWR VPWR VGND _1099_ _1098_ _1088_ _1095_ sky130_fd_sc_hd__mux2_1
X_7040_ VPWR VGND VPWR VGND _2138_ _3353_ _3352_ _2126_ _3354_ sky130_fd_sc_hd__or4_1
X_4183_ VPWR VGND _1030_ _1029_ VPWR VGND sky130_fd_sc_hd__buf_2
X_7942_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[1\] clknet_leaf_50_clk _0055_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7873_ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[28\] clknet_leaf_48_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[28\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6824_ VPWR VGND VGND VPWR _3195_ _3197_ _3196_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_159 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6755_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[21\] _3134_
+ net31 sky130_fd_sc_hd__nand2_1
X_3967_ VPWR VGND VGND VPWR _0817_ _0819_ _0818_ sky130_fd_sc_hd__nand2_1
X_5706_ VPWR VGND VPWR VGND _2358_ net188 sky130_fd_sc_hd__inv_2
XFILLER_0_73_641 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_70_72 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.i_regbuf\[27\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[27\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[31\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_343 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_30_clk VGND VPWR clknet_3_7__leaf_clk clknet_leaf_30_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_6686_ VGND VPWR VGND VPWR _0447_ _0883_ _3027_ _3071_ _2061_ sky130_fd_sc_hd__o211a_1
X_3898_ VPWR VGND VPWR VGND _0617_ _0749_ _0615_ _0750_ i_tinyqv.cpu.instr_data_start\[13\]
+ sky130_fd_sc_hd__a22o_1
X_8425_ i_tinyqv.cpu.i_core.imm_lo\[3\] clknet_leaf_23_clk _0523_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_2
X_5637_ VGND VPWR VPWR VGND _2311_ i_tinyqv.cpu.instr_data_in\[3\] _2309_ net260 sky130_fd_sc_hd__mux2_1
X_5568_ VGND VPWR _2259_ _2242_ _2261_ net142 VPWR VGND sky130_fd_sc_hd__o21ai_1
X_8356_ i_tinyqv.cpu.instr_data_start\[14\] clknet_leaf_36_clk _0455_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
Xhold141 net170 i_uart_tx.cycle_counter\[8\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_8287_ i_tinyqv.mem.qspi_data_buf\[27\] clknet_leaf_17_clk _0386_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_4519_ VPWR VGND VPWR VGND i_tinyqv.mem.data_from_read\[18\] _0689_ _1358_ _0748_
+ i_tinyqv.mem.data_from_read\[22\] _0957_ sky130_fd_sc_hd__a221o_1
Xhold152 net181 i_tinyqv.cpu.data_addr\[13\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7307_ VPWR VGND VPWR VGND _3438_ _0624_ _3579_ _0560_ sky130_fd_sc_hd__a21o_1
Xhold130 net159 i_tinyqv.cpu.i_core.mcause\[1\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 net214 i_uart_tx.cycle_counter\[6\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5499_ VGND VPWR _0121_ _2211_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7238_ VGND VPWR _0547_ _3523_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xhold174 net203 i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[25\] VPWR VGND VGND
+ VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 net192 i_tinyqv.cpu.i_core.mip\[17\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.i_regbuf\[16\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[16\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[20\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 net225 i_uart_rx.recieved_data\[2\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7169_ VPWR VGND VGND VPWR _3471_ _3446_ _3470_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_660 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_21_clk VGND VPWR clknet_3_3__leaf_clk clknet_leaf_21_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_0_51_368 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4870_ VGND VPWR VPWR VGND _1677_ i_tinyqv.cpu.debug_rd\[2\] _1674_ i_tinyqv.cpu.i_core.i_registers.reg_access\[8\]\[2\]
+ sky130_fd_sc_hd__mux2_1
X_3821_ VPWR VGND VPWR VGND _0669_ _0672_ _0665_ _0673_ sky130_fd_sc_hd__or3_1
X_6540_ VGND VPWR VPWR VGND _2951_ _2322_ _2925_ _2950_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_12_clk VGND VPWR clknet_3_2__leaf_clk clknet_leaf_12_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_0_15_505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_6471_ VGND VPWR VGND VPWR _2894_ _2625_ _2893_ _2647_ _0845_ sky130_fd_sc_hd__a211o_1
XFILLER_0_2_421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5422_ VPWR VGND VPWR VGND _2152_ _2149_ _2151_ sky130_fd_sc_hd__or2_2
X_8210_ i_tinyqv.cpu.i_core.i_shift.a\[31\] clknet_leaf_40_clk _0322_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
X_5353_ VPWR VGND VGND VPWR _2090_ i_tinyqv.cpu.i_core.mepc\[0\] net18 sky130_fd_sc_hd__or2_1
X_8141_ i_tinyqv.cpu.data_addr\[16\] clknet_leaf_34_clk _0253_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_4304_ VPWR VGND VPWR VGND _1120_ _1083_ _1150_ _1151_ sky130_fd_sc_hd__a21oi_1
X_5284_ VPWR VGND VPWR VGND _2008_ _2005_ _2034_ _2036_ sky130_fd_sc_hd__a21o_1
X_8072_ i_tinyqv.cpu.i_core.mie\[19\] clknet_leaf_37_clk _0207_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_4235_ VGND VPWR VPWR VGND _1082_ i_tinyqv.cpu.i_core.i_shift.a\[29\] _1036_ i_tinyqv.cpu.i_core.i_shift.a\[2\]
+ sky130_fd_sc_hd__mux2_1
X_7023_ VPWR VGND VGND VPWR _2067_ _3339_ _0516_ sky130_fd_sc_hd__nor2_1
X_4166_ VGND VPWR VPWR VGND _1013_ _1011_ _1012_ _0976_ sky130_fd_sc_hd__mux2_1
X_4097_ VPWR VGND VGND VPWR _0942_ _0916_ _0944_ _0933_ sky130_fd_sc_hd__nor3_4
X_7925_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[16\] clknet_leaf_36_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[16\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7856_ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[11\] clknet_leaf_45_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[11\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6807_ VGND VPWR VGND VPWR _3182_ _3040_ _3180_ _3181_ _3047_ sky130_fd_sc_hd__o211a_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.i_regbuf\[28\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[28\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_37_107 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4999_ VPWR VGND VGND VPWR _1763_ _1762_ _1760_ sky130_fd_sc_hd__or2_1
X_7787_ i_tinyqv.cpu.i_core.i_registers.reg_access\[7\]\[2\] clknet_leaf_52_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[6\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6738_ VGND VPWR _3118_ _3119_ _3116_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_6669_ VGND VPWR _3055_ _3056_ _3054_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_8408_ i_tinyqv.cpu.counter\[3\] clknet_leaf_24_clk _0506_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_33_357 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_8339_ i_tinyqv.mem.q_ctrl.addr\[1\] clknet_leaf_33_clk _0438_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.i_regbuf\[17\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[17\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[21\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.i_regbuf\[31\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[31\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[3\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.i_regbuf\[20\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[20\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[24\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_655 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.i_regbuf\[16\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[16\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[20\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_instrret.i_regbuf\[30\] i_tinyqv.cpu.i_core.i_instrret.reg_buf\[30\]
+ i_tinyqv.cpu.i_core.i_instrret.register\[2\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_cycles.i_regbuf\[14\] i_tinyqv.cpu.i_core.i_cycles.reg_buf\[14\]
+ i_tinyqv.cpu.i_core.i_cycles.register\[18\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4020_ VPWR VGND _0870_ _0869_ _0868_ VPWR VGND sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_1_clk VGND VPWR clknet_3_0__leaf_clk clknet_leaf_1_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_5971_ VGND VPWR VPWR VGND _2546_ i_tinyqv.cpu.i_core.mepc\[21\] _2107_ i_tinyqv.cpu.i_core.i_shift.a\[25\]
+ sky130_fd_sc_hd__mux2_1
X_4922_ VPWR VGND _1707_ i_tinyqv.mem.q_ctrl.fsm_state\[0\] VPWR VGND sky130_fd_sc_hd__buf_2
X_7710_ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[25\] clknet_leaf_56_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[25\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7641_ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[20\] clknet_leaf_56_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[20\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4853_ VGND VPWR _0032_ _1667_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4784_ VPWR VGND _1619_ _0748_ VPWR VGND sky130_fd_sc_hd__buf_2
X_7572_ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[15\] clknet_leaf_58_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[15\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_3804_ VGND VPWR i_tinyqv.cpu.alu_op\[1\] _0656_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_6523_ VGND VPWR _0420_ _2935_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6454_ VGND VPWR VGND VPWR _0406_ _2855_ _2857_ net289 _2305_ sky130_fd_sc_hd__a211o_1
X_5405_ VPWR VGND VGND VPWR _1452_ _1493_ _2135_ sky130_fd_sc_hd__nor2_1
X_6385_ VGND VPWR VPWR VGND _2824_ _2823_ _2797_ i_tinyqv.mem.q_ctrl.delay_cycles_cfg\[2\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_349 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_8124_ i_spi.data\[7\] clknet_leaf_18_clk _0236_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5336_ VGND VPWR _2077_ i_tinyqv.cpu.i_core.time_hi\[0\] i_tinyqv.cpu.i_core.time_hi\[1\]
+ _2074_ VPWR VGND sky130_fd_sc_hd__and3_1
X_8055_ i_spi.clock_count\[0\] clknet_leaf_27_clk _0190_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5267_ VGND VPWR VGND VPWR _2020_ _1996_ _1969_ _1995_ sky130_fd_sc_hd__a21bo_1
X_4218_ VGND VPWR VPWR VGND _1065_ i_tinyqv.cpu.i_core.i_shift.a\[19\] _1027_ i_tinyqv.cpu.i_core.i_shift.a\[12\]
+ sky130_fd_sc_hd__mux2_1
X_7006_ VGND VPWR VGND VPWR _3305_ _1492_ _1491_ _1452_ _3325_ sky130_fd_sc_hd__and4bb_1
X_5198_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[12\] _1953_ _1167_ sky130_fd_sc_hd__nand2_1
X_4149_ VGND VPWR _0996_ _0995_ _0984_ _0987_ VPWR VGND sky130_fd_sc_hd__and3_1
X_7908_ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[31\] clknet_leaf_48_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[31\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7839_ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[26\] clknet_leaf_3_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[26\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.i_regbuf\[21\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[21\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[25\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.i_regbuf\[28\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[28\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_71_205 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_25_600 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_4_549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_6170_ VGND VPWR _0337_ _2665_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5121_ VPWR VGND VGND VPWR _1879_ _1855_ _1878_ sky130_fd_sc_hd__or2_1
X_5052_ VPWR VGND _1813_ _1789_ VPWR VGND sky130_fd_sc_hd__buf_2
X_4003_ VPWR VGND VGND VPWR i_tinyqv.cpu.no_write_in_progress _0854_ i_tinyqv.cpu.is_store
+ sky130_fd_sc_hd__nand2_4
XFILLER_0_75_500 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5954_ VGND VPWR VPWR VGND _2535_ _2534_ _2524_ i_tinyqv.cpu.data_addr\[15\] sky130_fd_sc_hd__mux2_1
X_5885_ VGND VPWR _0230_ _2487_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4905_ VGND VPWR _0058_ _1697_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4836_ VGND VPWR _0041_ _1657_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7624_ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[3\] clknet_leaf_1_clk _0045_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7555_ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[30\] clknet_leaf_46_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[30\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_633 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6506_ VPWR VGND VPWR VGND _1711_ _2920_ _2782_ i_tinyqv.mem.q_ctrl.read_cycles_count\[0\]
+ sky130_fd_sc_hd__or3b_2
XFILLER_0_43_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4767_ VGND VPWR VPWR VGND _1602_ _0610_ _1599_ _0916_ _1601_ sky130_fd_sc_hd__o2bb2a_1
X_4698_ VGND VPWR VPWR VGND _1533_ _1517_ _1516_ _1480_ _1534_ sky130_fd_sc_hd__or4_4
X_7486_ VPWR VGND VGND VPWR _3239_ _3228_ _3725_ sky130_fd_sc_hd__nor2_1
X_6437_ VGND VPWR VPWR VGND _2869_ _2864_ _2787_ _2801_ _2868_ _2790_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_30_135 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6368_ VPWR VGND _2809_ _2788_ _2784_ i_tinyqv.mem.q_ctrl.delay_cycles_cfg\[0\] _2808_
+ VGND VPWR sky130_fd_sc_hd__a31o_1
X_5319_ VPWR VGND VPWR VGND _1401_ _2064_ _2065_ _2063_ sky130_fd_sc_hd__o21bai_1
X_8107_ i_tinyqv.cpu.instr_data\[0\]\[7\] clknet_leaf_10_clk _0219_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_6299_ VGND VPWR VPWR VGND _2759_ _1720_ _1552_ i_tinyqv.mem.qspi_data_buf\[14\]
+ sky130_fd_sc_hd__mux2_1
X_8038_ i_debug_uart_tx.data_to_send\[0\] clknet_leaf_29_clk _0173_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
Xhold89 net118 i_tinyqv.cpu.data_out\[25\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 net107 i_tinyqv.cpu.data_out\[24\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 net96 i_tinyqv.cpu.data_addr\[11\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_9 _2938_ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_0_61_293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_21_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.i_regbuf\[6\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[6\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[10\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_533 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5670_ i_debug_uart_tx.cycle_counter\[4\] i_debug_uart_tx.cycle_counter\[3\] _2331_
+ i_debug_uart_tx.cycle_counter\[1\] VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_4621_ VPWR VGND VGND VPWR _1457_ i_tinyqv.cpu.instr_data\[3\]\[2\] _1422_ sky130_fd_sc_hd__or2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.i_regbuf\[4\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[4\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[8\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_25_485 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4552_ VPWR VGND VPWR VGND _1388_ i_tinyqv.cpu.i_core.mem_op\[0\] sky130_fd_sc_hd__inv_2
X_7340_ VGND VPWR VGND VPWR _0567_ i_tinyqv.cpu.instr_len\[1\] _3282_ _3312_ _1753_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_13_658 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_4483_ VPWR VGND VGND VPWR _1320_ _1322_ _1321_ sky130_fd_sc_hd__nand2_1
X_7271_ VPWR VGND VPWR VGND _3548_ _3460_ _3532_ _3549_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_157 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6222_ VGND VPWR VPWR VGND _2700_ _2702_ _2701_ sky130_fd_sc_hd__xor2_1
XFILLER_0_21_680 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_585 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6153_ VGND VPWR VPWR VGND _2657_ i_tinyqv.cpu.i_core.mepc\[4\] _2656_ i_tinyqv.cpu.i_core.mepc\[0\]
+ sky130_fd_sc_hd__mux2_1
X_5104_ VPWR VGND VGND VPWR _1863_ i_tinyqv.cpu.i_core.multiplier.accum\[8\] _1861_
+ sky130_fd_sc_hd__or2_1
X_6084_ VGND VPWR VPWR VGND _2610_ i_tinyqv.cpu.i_core.i_shift.a\[14\] _2596_ i_tinyqv.cpu.i_core.i_shift.a\[18\]
+ sky130_fd_sc_hd__mux2_1
X_5035_ VGND VPWR _1796_ _1797_ i_tinyqv.cpu.i_core.multiplier.accum\[5\] VPWR VGND
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6986_ VPWR VGND VGND VPWR _3308_ _3307_ _1514_ sky130_fd_sc_hd__nor2b_2
X_5937_ VGND VPWR VPWR VGND _2523_ i_tinyqv.cpu.i_core.mepc\[10\] _2504_ i_tinyqv.cpu.i_core.i_shift.a\[14\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_641 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7607_ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[18\] clknet_leaf_2_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[18\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.i_regbuf\[10\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[10\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[14\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5868_ VGND VPWR _0222_ _2478_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5799_ VPWR VGND VPWR VGND _2427_ net162 _2429_ _0203_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_162 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_4819_ VPWR VGND _1189_ _1648_ _1647_ VPWR VGND sky130_fd_sc_hd__and2_2
X_7538_ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[13\] clknet_leaf_47_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[13\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7469_ VGND VPWR _2682_ _3005_ _3711_ net288 VPWR VGND sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_19_Right_19 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_39_533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_39_588 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_54_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_3_1__f_clk VGND VPWR VGND VPWR clknet_0_clk clknet_3_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_28_Right_28 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Right_37 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6840_ VGND VPWR VPWR VGND _3212_ _3211_ _2990_ _2544_ sky130_fd_sc_hd__mux2_1
X_6771_ _3149_ _3147_ _3148_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_5722_ VPWR VGND VGND VPWR _2370_ _2339_ _2333_ sky130_fd_sc_hd__or2_1
X_8510_ i_tinyqv.cpu.i_core.i_instrret.register\[16\] clknet_leaf_49_clk i_tinyqv.cpu.i_core.i_instrret.reg_buf\[16\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_3983_ VGND VPWR VGND VPWR _0835_ _0820_ _0834_ _0656_ net141 sky130_fd_sc_hd__a211o_1
X_5653_ VGND VPWR i_tinyqv.cpu.instr_data_in\[10\] _2320_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_8441_ i_tinyqv.cpu.imm\[19\] clknet_leaf_21_clk _0539_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_33_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5584_ VGND VPWR VGND VPWR _0147_ net240 _2263_ _2270_ _2240_ sky130_fd_sc_hd__o211a_1
X_8372_ i_tinyqv.cpu.data_continue clknet_leaf_21_clk _0028_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4604_ VGND VPWR VPWR VGND i_tinyqv.cpu.additional_mem_ops\[1\] i_tinyqv.cpu.additional_mem_ops\[0\]
+ i_tinyqv.cpu.additional_mem_ops\[2\] _1440_ sky130_fd_sc_hd__or3_2
XPHY_EDGE_ROW_46_Right_46 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4535_ VPWR VGND VGND VPWR _0907_ _1371_ _0909_ _1373_ _1374_ sky130_fd_sc_hd__o22a_1
X_7323_ VPWR VGND VPWR VGND _0711_ i_tinyqv.cpu.mem_op_increment_reg _3591_ _3592_
+ sky130_fd_sc_hd__a21oi_1
X_4466_ VPWR VGND uo_out[2] _1306_ VPWR VGND sky130_fd_sc_hd__buf_4
X_7254_ _3535_ _1507_ _3300_ _3314_ _2121_ VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_4397_ VPWR VGND VGND VPWR _0724_ _1235_ _1239_ _1240_ sky130_fd_sc_hd__o21a_1
X_6205_ VGND VPWR _0350_ _2687_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7185_ VPWR VGND VPWR VGND _3438_ net231 _3483_ _0534_ sky130_fd_sc_hd__a21o_1
X_6136_ VPWR VGND VPWR VGND _2642_ _2641_ _2643_ _2644_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_55_Right_55 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6067_ VGND VPWR _0298_ _2601_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5018_ VPWR VGND VGND VPWR _1570_ _1781_ _1577_ sky130_fd_sc_hd__nand2_1
X_6969_ VGND VPWR VGND VPWR _3292_ _2124_ _1473_ _1426_ _1420_ sky130_fd_sc_hd__and4_2
XPHY_EDGE_ROW_64_Right_64 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_23_219 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_73_Right_73 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_80_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.i_regbuf\[10\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[10\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[14\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_4320_ VGND VPWR _1166_ _1167_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_4251_ VGND VPWR VPWR VGND _1098_ _1097_ _1083_ _1096_ sky130_fd_sc_hd__mux2_1
X_4182_ VGND VPWR _1028_ _1029_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_7941_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[0\] clknet_leaf_50_clk _0054_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7872_ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[27\] clknet_leaf_48_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[27\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6823_ VPWR VGND VGND VPWR _3196_ i_tinyqv.cpu.instr_data_start\[19\] i_tinyqv.cpu.imm\[19\]
+ sky130_fd_sc_hd__or2_1
X_6754_ VGND VPWR VGND VPWR _0453_ _0726_ _3123_ _3133_ _3093_ sky130_fd_sc_hd__o211a_1
X_3966_ VPWR VGND VGND VPWR net86 _0818_ _0816_ sky130_fd_sc_hd__nand2_1
X_5705_ VGND VPWR VGND VPWR _0181_ i_debug_uart_tx.cycle_counter\[0\] _0989_ _2356_
+ _2357_ sky130_fd_sc_hd__o211a_1
X_6685_ VPWR VGND VGND VPWR _3037_ _3071_ _3070_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_3897_ VGND VPWR i_tinyqv.cpu.pc\[1\] _0749_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_5636_ VGND VPWR _0159_ _2310_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8424_ i_tinyqv.cpu.i_core.imm_lo\[2\] clknet_leaf_9_clk _0522_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_2
X_5567_ VPWR VGND VGND VPWR _2259_ _2260_ _0140_ sky130_fd_sc_hd__nor2_1
X_8355_ i_tinyqv.cpu.instr_data_start\[13\] clknet_leaf_36_clk _0454_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_13_241 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold131 net160 i_uart_rx.recieved_data\[5\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 net171 _2219_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5498_ _2209_ _2199_ _2211_ _2210_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
Xhold120 net149 i_tinyqv.cpu.data_out\[12\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_8286_ i_tinyqv.mem.qspi_data_buf\[26\] clknet_leaf_14_clk _0385_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_7306_ VGND VPWR VGND VPWR _3579_ _2140_ _3491_ _3578_ _3359_ sky130_fd_sc_hd__o211a_1
X_4518_ VPWR VGND VPWR VGND _1347_ _0814_ _0880_ _1357_ _1356_ sky130_fd_sc_hd__a22o_1
Xhold153 net182 i_tinyqv.cpu.i_core.mie\[17\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 net193 i_uart_rx.rxd_reg\[1\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 net204 i_spi.clock_divider\[1\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7237_ VGND VPWR VPWR VGND _3523_ _3522_ _3396_ i_tinyqv.cpu.imm\[27\] sky130_fd_sc_hd__mux2_1
Xhold186 net215 i_tinyqv.cpu.i_core.i_registers.reg_access\[12\]\[0\] VPWR VGND VGND
+ VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4449_ VGND VPWR VPWR VGND _1292_ _1145_ _1088_ _1131_ sky130_fd_sc_hd__mux2_1
Xhold197 net226 i_tinyqv.cpu.i_core.mepc\[13\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7168_ VGND VPWR VPWR VGND _3469_ _3447_ _3445_ _3470_ sky130_fd_sc_hd__or3b_1
X_6119_ VPWR VGND VPWR VGND i_tinyqv.cpu.i_core.i_shift.a\[30\] _2596_ _0321_ _2628_
+ _2629_ _2630_ sky130_fd_sc_hd__a221o_1
X_7099_ VPWR VGND VGND VPWR _3368_ i_tinyqv.cpu.instr_data\[1\]\[8\] _3366_ i_tinyqv.cpu.instr_data\[0\]\[8\]
+ _3408_ _3407_ sky130_fd_sc_hd__o221a_1
XFILLER_0_49_683 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_48_182 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_17_591 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_66 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_3820_ VGND VPWR VPWR VGND _0672_ _0670_ _0667_ i_tinyqv.cpu.i_core.i_registers.reg_access\[2\]\[3\]
+ net25 i_tinyqv.cpu.i_core.i_registers.reg_access\[8\]\[3\] sky130_fd_sc_hd__a32o_1
XFILLER_0_55_631 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_70_612 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_40_32 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_70_645 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6470_ VPWR VGND VGND VPWR _1260_ _2625_ _2893_ sky130_fd_sc_hd__nor2_1
X_5421_ VPWR VGND VGND VPWR _1399_ _1443_ _2150_ _2151_ sky130_fd_sc_hd__o21a_1
X_8140_ i_tinyqv.cpu.data_addr\[15\] clknet_leaf_34_clk _0252_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_5352_ VPWR VGND VGND VPWR _2088_ _0922_ _0937_ _2089_ sky130_fd_sc_hd__nor3_1
X_4303_ VPWR VGND VGND VPWR _1083_ _1086_ _1150_ sky130_fd_sc_hd__nor2_1
X_8071_ i_tinyqv.cpu.i_core.mip\[16\] clknet_leaf_23_clk _0206_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_5283_ VPWR VGND VGND VPWR _2005_ _2008_ _2035_ _2034_ sky130_fd_sc_hd__nand3_1
X_7022_ VPWR VGND VPWR VGND _3335_ _3333_ _3338_ _3339_ sky130_fd_sc_hd__a21oi_1
X_4234_ VGND VPWR VPWR VGND _1081_ i_tinyqv.cpu.i_core.i_shift.a\[28\] _1029_ i_tinyqv.cpu.i_core.i_shift.a\[3\]
+ sky130_fd_sc_hd__mux2_1
X_4165_ VPWR VGND VGND VPWR _1012_ _0869_ _0979_ sky130_fd_sc_hd__nand2_2
XFILLER_0_65_73 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4096_ VPWR VGND VGND VPWR _0942_ _0937_ _0916_ _0943_ sky130_fd_sc_hd__nor3_1
X_7924_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[15\] clknet_leaf_24_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[15\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7855_ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[10\] clknet_leaf_5_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[10\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6806_ VPWR VGND VGND VPWR _1390_ _3181_ _2538_ sky130_fd_sc_hd__nand2_1
X_4998_ VPWR VGND _1762_ _1761_ i_tinyqv.cpu.is_store VPWR VGND sky130_fd_sc_hd__and2_1
X_7786_ i_tinyqv.cpu.i_core.i_registers.reg_access\[7\]\[1\] clknet_leaf_52_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[5\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6737_ VPWR VGND VGND VPWR _3105_ _3117_ _3118_ sky130_fd_sc_hd__nor2_1
X_3949_ VPWR VGND VPWR VGND i_tinyqv.cpu.i_core.i_registers.reg_access\[15\]\[2\]
+ _0677_ _0801_ _0684_ i_tinyqv.cpu.i_core.i_registers.reg_access\[13\]\[2\] _0800_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6668_ VPWR VGND VGND VPWR _3043_ _3044_ _3041_ _3055_ sky130_fd_sc_hd__o21a_1
X_5619_ VPWR VGND VGND VPWR _2298_ i_uart_rx.fsm_state\[3\] _2281_ sky130_fd_sc_hd__or2_1
X_6599_ VPWR VGND VGND VPWR _2994_ _2996_ _2061_ _0435_ sky130_fd_sc_hd__o21a_1
X_8407_ i_tinyqv.cpu.counter\[2\] clknet_leaf_22_clk _0505_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_8338_ i_tinyqv.mem.q_ctrl.addr\[0\] clknet_leaf_29_clk _0437_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_8269_ i_tinyqv.mem.qspi_data_buf\[9\] clknet_leaf_14_clk _0368_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.i_regbuf\[24\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[24\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[28\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.i_regbuf\[13\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[13\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[17\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_49_480 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_52_689 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xi_tinyqv.cpu.i_core.i_instrret.i_regbuf\[23\] i_tinyqv.cpu.i_core.i_instrret.reg_buf\[23\]
+ i_tinyqv.cpu.i_core.i_instrret.register\[27\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5970_ VGND VPWR _0257_ _2545_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4921_ VGND VPWR i_tinyqv.mem.q_ctrl.fsm_state\[2\] _1706_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_4852_ VGND VPWR VPWR VGND _1667_ i_tinyqv.cpu.debug_rd\[2\] _1664_ i_tinyqv.cpu.i_core.i_registers.reg_access\[10\]\[2\]
+ sky130_fd_sc_hd__mux2_1
X_7640_ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[19\] clknet_leaf_46_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[19\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_3803_ VGND VPWR VPWR VGND _0655_ _0654_ _0652_ _0623_ sky130_fd_sc_hd__mux2_4
X_4783_ VGND VPWR VGND VPWR _1618_ uo_out[7] _1617_ _1001_ _0971_ sky130_fd_sc_hd__a211o_1
XFILLER_0_55_461 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_7571_ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[14\] clknet_leaf_54_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[14\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_6522_ VGND VPWR VPWR VGND _2935_ _2318_ _2925_ _2934_ sky130_fd_sc_hd__mux2_1
X_6453_ VPWR VGND VPWR VGND _2838_ _2840_ _0405_ _2855_ net208 _2305_ sky130_fd_sc_hd__a221o_1
X_5404_ VPWR VGND VPWR VGND _2130_ _2133_ _2131_ _2126_ _2134_ sky130_fd_sc_hd__or4_1
XFILLER_0_42_177 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6384_ VPWR VGND VGND VPWR i_tinyqv.mem.q_ctrl.read_cycles_count\[0\] i_tinyqv.mem.q_ctrl.read_cycles_count\[1\]
+ i_tinyqv.mem.q_ctrl.read_cycles_count\[2\] _2823_ sky130_fd_sc_hd__o21a_1
X_8123_ i_spi.data\[6\] clknet_leaf_18_clk _0235_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_564 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_5335_ VPWR VGND VGND VPWR _2075_ _2076_ _0092_ sky130_fd_sc_hd__nor2_1
X_8054_ i_debug_uart_tx.fsm_state\[3\] clknet_leaf_30_clk _0189_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5266_ VPWR VGND _2019_ _2018_ _2017_ VPWR VGND sky130_fd_sc_hd__and2_1
X_4217_ VGND VPWR VPWR VGND _1064_ i_tinyqv.cpu.i_core.i_shift.a\[18\] _1027_ i_tinyqv.cpu.i_core.i_shift.a\[13\]
+ sky130_fd_sc_hd__mux2_1
X_7005_ VGND VPWR VGND VPWR _0513_ _3312_ _3320_ _3324_ _3205_ sky130_fd_sc_hd__o211a_1
X_5197_ VGND VPWR _1951_ _1952_ _1950_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_4148_ VPWR VGND VPWR VGND _0995_ _0969_ sky130_fd_sc_hd__inv_2
X_4079_ VPWR VGND VPWR VGND _0923_ _0925_ _0924_ i_tinyqv.cpu.i_core.imm_lo\[6\] _0926_
+ sky130_fd_sc_hd__or4_1
X_7907_ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[30\] clknet_leaf_2_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[30\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7838_ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[25\] clknet_leaf_3_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[25\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7769_ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[20\] clknet_leaf_0_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[20\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.i_regbuf\[25\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[25\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[29\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.i_regbuf\[14\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[14\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[18\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_612 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_24_122 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_52_464 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_5120_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[7\] _1878_ _1789_ sky130_fd_sc_hd__nand2_1
X_5051_ VGND VPWR VPWR VGND _1810_ _1812_ _1811_ sky130_fd_sc_hd__xor2_1
X_4002_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.is_interrupt i_tinyqv.cpu.is_branch
+ _0853_ sky130_fd_sc_hd__nor2_1
X_5953_ VGND VPWR VPWR VGND _2534_ i_tinyqv.cpu.i_core.mepc\[15\] _2107_ i_tinyqv.cpu.i_core.i_shift.a\[19\]
+ sky130_fd_sc_hd__mux2_1
X_5884_ VGND VPWR VPWR VGND _2487_ _2486_ _2399_ i_spi.data\[1\] sky130_fd_sc_hd__mux2_1
XFILLER_0_62_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4904_ VGND VPWR VPWR VGND _1697_ _1184_ _1696_ i_tinyqv.cpu.i_core.i_registers.reg_access\[2\]\[0\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_47_236 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4835_ VGND VPWR VPWR VGND _1657_ net32 _1653_ net101 sky130_fd_sc_hd__mux2_1
XFILLER_0_7_333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7623_ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[2\] clknet_leaf_1_clk _0044_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_355 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_7554_ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[29\] clknet_leaf_54_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[29\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4766_ VPWR VGND VGND VPWR _1601_ _0899_ _1600_ sky130_fd_sc_hd__or2_1
X_6505_ VGND VPWR VPWR VGND _2919_ i_tinyqv.mem.q_ctrl.spi_in_buffer\[0\] _2918_ i_tinyqv.mem.q_ctrl.spi_in_buffer\[4\]
+ sky130_fd_sc_hd__mux2_1
X_7485_ VPWR VGND VGND VPWR _3723_ _2733_ _3625_ i_tinyqv.mem.q_ctrl.addr\[21\] _0593_
+ _3724_ sky130_fd_sc_hd__o221a_1
X_4697_ VPWR VGND _1533_ _1532_ i_tinyqv.cpu.instr_fetch_started VPWR VGND sky130_fd_sc_hd__and2_1
X_6436_ VPWR VGND VPWR VGND _1708_ _1714_ _2867_ _2868_ sky130_fd_sc_hd__a21oi_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.i_regbuf\[7\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[7\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[11\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_6367_ VGND VPWR _2801_ _2804_ _2799_ _2808_ _2807_ _2787_ VPWR VGND sky130_fd_sc_hd__a41o_1
X_8106_ i_tinyqv.cpu.instr_data\[0\]\[6\] clknet_leaf_4_clk _0218_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5318_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.is_interrupt _2064_ _0744_ sky130_fd_sc_hd__nand2_1
X_6298_ VGND VPWR _0372_ _2758_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8037_ i_tinyqv.cpu.instr_data\[3\]\[15\] clknet_leaf_12_clk _0172_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5249_ VGND VPWR VPWR VGND _2000_ _2002_ _2001_ sky130_fd_sc_hd__xor2_1
Xhold68 VGND VPWR i_debug_uart_tx.uart_tx_data\[1\] net97 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xhold79 net108 i_tinyqv.cpu.i_core.time_hi\[2\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_247 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.i_regbuf\[6\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[6\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[10\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4620_ VPWR VGND VGND VPWR _1452_ _1456_ _1455_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_325 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4551_ VPWR VGND VGND VPWR _1386_ _1387_ _0908_ sky130_fd_sc_hd__nor2_2
XFILLER_0_12_136 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4482_ VGND VPWR _1251_ _1247_ _1321_ _1249_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_7270_ VPWR VGND VPWR VGND _3299_ _1473_ _3304_ _3548_ sky130_fd_sc_hd__a21o_1
X_6221_ VPWR VGND VGND VPWR _1060_ _2701_ _1845_ sky130_fd_sc_hd__nand2_1
X_6152_ VPWR VGND _2656_ _1386_ VPWR VGND sky130_fd_sc_hd__buf_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.i_regbuf\[4\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[4\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[8\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5103_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.multiplier.accum\[8\] _1862_ _1861_
+ sky130_fd_sc_hd__nand2_1
X_6083_ VGND VPWR _0306_ _2609_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5034_ VGND VPWR VPWR VGND _1793_ _1796_ _1795_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_69_Left_150 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6985_ VPWR VGND VGND VPWR _3307_ _1502_ _1510_ sky130_fd_sc_hd__or2_1
X_5936_ VGND VPWR _0246_ _2522_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7606_ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[17\] clknet_leaf_52_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[17\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_206 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5867_ VGND VPWR VPWR VGND _2478_ i_tinyqv.cpu.instr_data\[0\]\[10\] _2469_ _2320_
+ sky130_fd_sc_hd__mux2_1
X_5798_ VPWR VGND _2429_ _1725_ _1004_ i_debug_uart_tx.uart_tx_data\[0\] _2229_ VGND
+ VPWR sky130_fd_sc_hd__a31o_1
X_4818_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_registers.rd\[1\] _1640_ _1647_
+ sky130_fd_sc_hd__nor2_1
X_7537_ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[12\] clknet_leaf_47_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[12\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4749_ VGND VPWR VPWR VGND _1322_ _1584_ net82 sky130_fd_sc_hd__xor2_1
X_7468_ VGND VPWR VGND VPWR _3710_ _3239_ _3199_ _3709_ _2682_ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6419_ VGND VPWR VGND VPWR _2854_ _2852_ _2853_ _1540_ _2844_ sky130_fd_sc_hd__a211o_1
X_7399_ VPWR VGND VGND VPWR _3017_ _3651_ _3652_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_618 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6770_ VPWR VGND VGND VPWR i_tinyqv.cpu.instr_data_start\[14\] _3148_ i_tinyqv.cpu.imm\[14\]
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_417 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_3982_ VPWR VGND VPWR VGND _0833_ _0832_ _0656_ _0834_ sky130_fd_sc_hd__a21oi_1
X_5721_ VPWR VGND VPWR VGND _2368_ _0988_ _2341_ _2369_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_76 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_8440_ i_tinyqv.cpu.imm\[18\] clknet_leaf_22_clk _0538_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_5652_ VGND VPWR _0166_ _2319_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5583_ VPWR VGND VGND VPWR _2270_ i_uart_rx.recieved_data\[5\] _2264_ sky130_fd_sc_hd__or2_1
X_8371_ i_tinyqv.cpu.data_read_n\[1\] clknet_leaf_20_clk _0470_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_4603_ VPWR VGND VGND VPWR _0837_ _1439_ _0863_ sky130_fd_sc_hd__nand2_1
X_4534_ VGND VPWR VPWR VGND _1373_ _1372_ _1012_ _1360_ sky130_fd_sc_hd__mux2_1
X_7322_ VPWR VGND VPWR VGND i_tinyqv.cpu.mem_op_increment_reg _0662_ _0663_ _3591_
+ sky130_fd_sc_hd__a21oi_1
X_4465_ VGND VPWR VPWR VGND _1306_ gpio_out\[2\] gpio_out_sel\[2\] _1305_ sky130_fd_sc_hd__mux2_1
X_7253_ VPWR VGND VPWR VGND _3533_ _2123_ _3335_ _3534_ _3299_ sky130_fd_sc_hd__a22o_1
X_4396_ VPWR VGND VGND VPWR _0909_ _1237_ _0907_ _1238_ _1239_ sky130_fd_sc_hd__o22a_1
X_6204_ VGND VPWR VPWR VGND _2687_ _2683_ _2686_ _1635_ sky130_fd_sc_hd__mux2_1
X_7184_ VGND VPWR _3483_ _3480_ _3359_ _3482_ VPWR VGND sky130_fd_sc_hd__and3_1
X_6135_ VPWR VGND VGND VPWR _0707_ _2642_ _2643_ sky130_fd_sc_hd__nor2_1
X_6066_ VGND VPWR VPWR VGND _2601_ i_tinyqv.cpu.i_core.i_shift.a\[9\] _2593_ i_tinyqv.cpu.i_core.i_shift.a\[5\]
+ sky130_fd_sc_hd__mux2_1
X_5017_ VPWR VGND _1780_ _1779_ _1778_ VPWR VGND sky130_fd_sc_hd__xor2_2
X_6968_ VGND VPWR _3290_ _3291_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_6899_ VPWR VGND VPWR VGND _3257_ net16 sky130_fd_sc_hd__inv_2
X_5919_ VGND VPWR VPWR VGND _2511_ i_tinyqv.cpu.i_core.mepc\[4\] _2504_ i_tinyqv.cpu.i_core.i_shift.a\[8\]
+ sky130_fd_sc_hd__mux2_1
X_8569_ VGND VPWR uio_oe[5] uio_oe[4] VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_32_710 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_16_261 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_16_272 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_7_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_2_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_22_231 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4250_ VGND VPWR VPWR VGND _1097_ i_tinyqv.cpu.i_core.i_shift.a\[27\] _1029_ i_tinyqv.cpu.i_core.i_shift.a\[4\]
+ sky130_fd_sc_hd__mux2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.i_regbuf\[28\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[28\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4181_ VGND VPWR _1027_ _1028_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_7940_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[31\] clknet_leaf_49_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[31\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7871_ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[26\] clknet_leaf_3_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[26\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6822_ VPWR VGND VGND VPWR i_tinyqv.cpu.instr_data_start\[19\] _3195_ i_tinyqv.cpu.imm\[19\]
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6753_ VPWR VGND VGND VPWR _3037_ _3133_ _3132_ sky130_fd_sc_hd__nand2_1
X_3965_ VPWR VGND VGND VPWR _0817_ net86 _0816_ sky130_fd_sc_hd__or2_1
X_5704_ VPWR VGND VGND VPWR _2198_ _2333_ _2357_ sky130_fd_sc_hd__nor2_1
X_6684_ VPWR VGND VPWR VGND _3062_ _3039_ _3070_ _2995_ _1340_ _3069_ sky130_fd_sc_hd__a221o_1
X_3896_ VPWR VGND _0748_ _0619_ VPWR VGND sky130_fd_sc_hd__buf_4
X_5635_ VGND VPWR VPWR VGND _2310_ i_tinyqv.cpu.instr_data_in\[2\] _2309_ net263 sky130_fd_sc_hd__mux2_1
X_8423_ i_tinyqv.cpu.i_core.imm_lo\[1\] clknet_leaf_7_clk _0521_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_2
X_5566_ VGND VPWR _2256_ _2242_ _2260_ net247 VPWR VGND sky130_fd_sc_hd__o21ai_1
X_8354_ i_tinyqv.cpu.instr_data_start\[12\] clknet_leaf_36_clk _0453_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
Xhold110 net139 _0084_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 net172 i_uart_rx.recieved_data\[7\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5497_ VPWR VGND _2210_ _2203_ i_uart_tx.cycle_counter\[3\] i_uart_tx.cycle_counter\[4\]
+ i_uart_tx.cycle_counter\[5\] VGND VPWR sky130_fd_sc_hd__a31o_1
X_8285_ i_tinyqv.mem.qspi_data_buf\[25\] clknet_leaf_14_clk _0384_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
Xhold132 net161 i_tinyqv.cpu.data_addr\[17\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_275 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold121 net150 i_tinyqv.cpu.i_core.i_registers.reg_access\[7\]\[2\] VPWR VGND VGND
+ VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7305_ VGND VPWR VGND VPWR _3578_ _3572_ _3573_ _1514_ _3577_ sky130_fd_sc_hd__a211o_1
X_4517_ VPWR VGND VPWR VGND _1355_ _0921_ _0880_ _1356_ sky130_fd_sc_hd__a21oi_1
Xhold176 net205 i_debug_uart_tx.data_to_send\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 net194 i_spi.bits_remaining\[3\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 net183 i_tinyqv.cpu.instr_fetch_started VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4448_ VPWR VGND VGND VPWR _1080_ _1291_ _1290_ sky130_fd_sc_hd__nand2_1
X_7236_ VPWR VGND _3522_ _3434_ _3330_ _3291_ _3510_ VGND VPWR sky130_fd_sc_hd__a31o_1
Xhold198 net227 i_tinyqv.cpu.imm\[15\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 net216 i_tinyqv.cpu.i_core.i_registers.reg_access\[7\]\[1\] VPWR VGND VGND
+ VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4379_ VGND VPWR VPWR VGND _1222_ _1221_ _0979_ _1220_ sky130_fd_sc_hd__mux2_1
X_7167_ VPWR VGND VGND VPWR _1478_ _2143_ _3298_ _3469_ sky130_fd_sc_hd__o21a_1
X_7098_ VPWR VGND VPWR VGND i_tinyqv.cpu.instr_data\[3\]\[8\] _3369_ _3407_ _3370_
+ i_tinyqv.cpu.instr_data\[2\]\[8\] _3372_ sky130_fd_sc_hd__a221o_1
X_6118_ _2630_ _1394_ i_tinyqv.cpu.i_core.mstatus_mte _0744_ _1392_ VGND VPWR VPWR
+ VGND sky130_fd_sc_hd__and4_1
X_6049_ VGND VPWR _0291_ _2590_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_610 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_55_643 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_39_194 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_54_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5420_ VPWR VGND VGND VPWR _1405_ _1438_ _2150_ sky130_fd_sc_hd__nor2_1
X_5351_ VPWR VGND VPWR VGND _2088_ _1124_ _0855_ sky130_fd_sc_hd__or2_2
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.i_regbuf\[29\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[29\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[1\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5282_ VPWR VGND VGND VPWR _2034_ _2032_ _2033_ sky130_fd_sc_hd__or2_1
X_4302_ VGND VPWR _1108_ _1149_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_8070_ i_tinyqv.cpu.i_core.mip\[17\] clknet_leaf_23_clk _0205_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_4233_ VPWR VGND _1080_ _1058_ VPWR VGND sky130_fd_sc_hd__buf_2
X_7021_ VGND VPWR VPWR VGND _3338_ _3337_ _3281_ i_tinyqv.cpu.is_branch sky130_fd_sc_hd__mux2_1
X_4164_ VGND VPWR VPWR VGND _1011_ i_tinyqv.cpu.instr_data_in\[4\] _0974_ i_tinyqv.cpu.instr_data_in\[0\]
+ sky130_fd_sc_hd__mux2_1
X_4095_ VGND VPWR VGND VPWR _0942_ i_tinyqv.cpu.i_core.imm_lo\[2\] i_tinyqv.cpu.i_core.imm_lo\[0\]
+ i_tinyqv.cpu.i_core.imm_lo\[1\] i_tinyqv.cpu.i_core.imm_lo\[3\] sky130_fd_sc_hd__or4b_4
X_7923_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[14\] clknet_leaf_25_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[14\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_201 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_7854_ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[9\] clknet_leaf_47_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[9\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6805_ VGND VPWR _3179_ _3180_ _3177_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_7785_ i_tinyqv.cpu.i_core.i_registers.reg_access\[7\]\[0\] clknet_leaf_1_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[4\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6736_ VGND VPWR VGND VPWR _3117_ _3095_ _3098_ _3106_ _3096_ sky130_fd_sc_hd__o211a_1
X_4997_ VPWR VGND VGND VPWR _1756_ _1761_ _0836_ sky130_fd_sc_hd__nor2_2
X_3948_ VPWR VGND VPWR VGND _0678_ i_tinyqv.cpu.i_core.i_registers.reg_access\[12\]\[2\]
+ _0674_ _0800_ i_tinyqv.cpu.i_core.i_registers.reg_access\[7\]\[2\] sky130_fd_sc_hd__a22o_1
X_6667_ VPWR VGND VGND VPWR _3052_ _3053_ _3054_ sky130_fd_sc_hd__nor2_1
X_3879_ VPWR VGND VPWR VGND _0646_ i_tinyqv.cpu.i_core.i_registers.reg_access\[13\]\[0\]
+ _0628_ _0731_ i_tinyqv.cpu.i_core.i_registers.reg_access\[10\]\[0\] sky130_fd_sc_hd__a22o_1
XFILLER_0_18_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_33_337 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5618_ VPWR VGND VPWR VGND _2296_ _2238_ _2280_ _2297_ sky130_fd_sc_hd__a21oi_1
X_8406_ i_tinyqv.cpu.data_out\[31\] clknet_leaf_20_clk _0504_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_6598_ _2996_ _1521_ _2995_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_5549_ VGND VPWR _0134_ _2248_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8337_ i_tinyqv.cpu.instr_write_offset\[2\] clknet_leaf_22_clk _0436_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.i_regbuf\[21\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[21\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[25\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_8268_ i_tinyqv.mem.qspi_data_buf\[8\] clknet_leaf_14_clk _0367_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_8199_ i_tinyqv.cpu.i_core.i_shift.a\[18\] clknet_leaf_40_clk _0311_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_7219_ VPWR VGND VGND VPWR _3511_ _3474_ i_tinyqv.cpu.imm\[20\] _3510_ _0540_ sky130_fd_sc_hd__o22a_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.i_regbuf\[17\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[17\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[21\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_37_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_36_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_23_Left_104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_19_89 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_instrret.i_regbuf\[16\] i_tinyqv.cpu.i_core.i_instrret.reg_buf\[16\]
+ i_tinyqv.cpu.i_core.i_instrret.register\[20\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_32_Left_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4920_ VGND VPWR _0057_ _1705_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_21 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_4851_ VGND VPWR _0031_ _1666_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_3802_ VGND VPWR VPWR VGND _0653_ _0654_ i_tinyqv.cpu.is_jal i_tinyqv.cpu.is_auipc
+ sky130_fd_sc_hd__o21ai_4
X_4782_ VPWR VGND VPWR VGND i_uart_rx.recieved_data\[7\] _0997_ _1617_ net14 gpio_out_sel\[7\]
+ _1616_ sky130_fd_sc_hd__a221o_1
X_7570_ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[13\] clknet_leaf_58_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[13\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6521_ VGND VPWR VPWR VGND _2934_ _2933_ _2792_ _2931_ sky130_fd_sc_hd__mux2_1
X_6452_ VPWR VGND VPWR VGND _2855_ net210 _2880_ _0404_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_41_Left_122 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5403_ VPWR VGND _2133_ _2132_ _2124_ VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_42_167 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6383_ VGND VPWR _0393_ _2822_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8122_ i_spi.data\[5\] clknet_leaf_18_clk _0234_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5334_ VGND VPWR _2074_ _2049_ _2076_ net246 VPWR VGND sky130_fd_sc_hd__o21ai_1
X_8053_ i_debug_uart_tx.fsm_state\[2\] clknet_leaf_30_clk _0188_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_5265_ VPWR VGND VGND VPWR _2018_ _2015_ _2016_ sky130_fd_sc_hd__or2_1
X_5196_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[10\] _1951_ _1880_ sky130_fd_sc_hd__nand2_1
X_4216_ VGND VPWR VPWR VGND _1063_ _1062_ _1050_ _1061_ sky130_fd_sc_hd__mux2_1
X_7004_ VGND VPWR VPWR VGND _3324_ _3323_ _3281_ i_tinyqv.cpu.is_store sky130_fd_sc_hd__mux2_1
X_4147_ VPWR VGND VPWR VGND net2 _0986_ _0994_ _0987_ _0993_ _0974_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_50_Left_131 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4078_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.imm_lo\[11\] _0925_ i_tinyqv.cpu.i_core.imm_lo\[10\]
+ sky130_fd_sc_hd__nand2_1
X_7906_ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[29\] clknet_leaf_2_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[29\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7837_ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[24\] clknet_leaf_48_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[24\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7768_ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[19\] clknet_leaf_58_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[19\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_462 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_6719_ VPWR VGND VGND VPWR _3102_ _3029_ _3101_ sky130_fd_sc_hd__or2_1
X_7699_ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[14\] clknet_leaf_53_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[14\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.i_regbuf\[22\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[22\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[26\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.i_regbuf\[29\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[29\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[1\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.i_regbuf\[18\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[18\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[22\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_101 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_4_529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.i_regbuf\[21\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[21\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[25\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5050_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[6\] _1811_ _1166_ sky130_fd_sc_hd__nand2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.i_regbuf\[10\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[10\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[14\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4001_ VPWR VGND VGND VPWR i_tinyqv.cpu.debug_instr_valid _0852_ i_tinyqv.cpu.is_auipc
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_20 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5952_ VGND VPWR _0251_ _2533_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4903_ _1641_ _1696_ _1188_ _1695_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_5883_ VGND VPWR VPWR VGND _2486_ i_spi.data\[0\] _2386_ i_debug_uart_tx.uart_tx_data\[1\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_97 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.i_regbuf\[9\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[9\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[13\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_708 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4834_ VGND VPWR _0040_ _1656_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7622_ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[1\] clknet_leaf_56_clk _0043_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4765_ VPWR VGND VPWR VGND _0898_ _0784_ i_tinyqv.cpu.instr_data_start\[19\] _1600_
+ sky130_fd_sc_hd__a21oi_1
X_7553_ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[28\] clknet_leaf_47_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[28\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6504_ VGND VPWR VGND VPWR i_tinyqv.mem.q_ctrl.read_cycles_count\[2\] i_tinyqv.mem.q_ctrl.read_cycles_count\[0\]
+ _2918_ _2789_ i_tinyqv.mem.q_ctrl.read_cycles_count\[1\] sky130_fd_sc_hd__or4bb_4
X_7484_ VPWR VGND VGND VPWR _3724_ i_tinyqv.mem.q_ctrl.addr\[17\] _3624_ sky130_fd_sc_hd__or2_1
X_4696_ VGND VPWR VGND VPWR _1532_ _1531_ i_tinyqv.mem.q_ctrl.data_ready _1530_ _0978_
+ sky130_fd_sc_hd__or4b_4
X_6435_ VPWR VGND VGND VPWR i_tinyqv.mem.q_ctrl.spi_flash_select _1713_ _1709_ _2867_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_551 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_3_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_6366_ VPWR VGND VPWR VGND _2806_ _2805_ i_tinyqv.mem.q_ctrl.read_cycles_count\[0\]
+ _2807_ sky130_fd_sc_hd__a21oi_1
X_8105_ i_tinyqv.cpu.instr_data\[0\]\[5\] clknet_leaf_3_clk _0217_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5317_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.mie\[18\] _2063_ _1228_ sky130_fd_sc_hd__nand2_1
X_6297_ VGND VPWR VPWR VGND _2758_ _1717_ _1552_ i_tinyqv.mem.qspi_data_buf\[13\]
+ sky130_fd_sc_hd__mux2_1
X_8036_ i_tinyqv.cpu.instr_data\[3\]\[14\] clknet_leaf_11_clk _0171_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5248_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[14\] _2001_ _1167_ sky130_fd_sc_hd__nand2_1
Xhold69 VGND VPWR i_debug_uart_tx.uart_tx_data\[2\] net98 VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_5179_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.multiplier.accum\[11\] _1935_ _1934_
+ sky130_fd_sc_hd__nand2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.i_regbuf\[7\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[7\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[11\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_7_Left_88 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_46_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_34_454 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_57_513 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_29_204 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_32_67 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_32_78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_65_590 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_25_443 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4550_ VPWR VGND VGND VPWR _1386_ _0688_ _0907_ sky130_fd_sc_hd__nand2_2
XFILLER_0_13_605 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_13_627 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_4481_ VGND VPWR VPWR VGND _1318_ _1320_ _1319_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_521 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_6220_ VPWR VGND VGND VPWR _2698_ _2700_ _2699_ sky130_fd_sc_hd__nand2_1
X_6151_ VGND VPWR _0328_ _2655_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5102_ VGND VPWR VPWR VGND _1859_ _1861_ _1860_ sky130_fd_sc_hd__xor2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.i_regbuf\[11\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[11\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[15\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6082_ VGND VPWR VPWR VGND _2609_ i_tinyqv.cpu.i_core.i_shift.a\[17\] _2592_ i_tinyqv.cpu.i_core.i_shift.a\[13\]
+ sky130_fd_sc_hd__mux2_1
X_5033_ VPWR VGND VPWR VGND _1768_ _1767_ _1794_ _1795_ sky130_fd_sc_hd__a21o_1
X_6984_ VPWR VGND VPWR VGND _1465_ _1492_ _2140_ _3306_ sky130_fd_sc_hd__or3_1
X_5935_ VGND VPWR VPWR VGND _2522_ _2521_ _2502_ i_tinyqv.cpu.data_addr\[9\] sky130_fd_sc_hd__mux2_1
X_5866_ VGND VPWR _0221_ _2477_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4817_ VGND VPWR _0049_ _1646_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7605_ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[16\] clknet_leaf_0_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[16\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5797_ VGND VPWR VGND VPWR _0202_ net98 _2427_ _2428_ _2221_ sky130_fd_sc_hd__o211a_1
XFILLER_0_8_687 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7536_ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[11\] clknet_leaf_45_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[11\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4748_ VGND VPWR VPWR VGND _1580_ _1583_ _1582_ sky130_fd_sc_hd__xor2_1
X_7467_ VPWR VGND VPWR VGND _3707_ _3708_ _3632_ _3709_ sky130_fd_sc_hd__or3_1
X_4679_ VGND VPWR VPWR VGND _1514_ _1511_ _1502_ _1495_ _1515_ sky130_fd_sc_hd__or4_4
X_6418_ VGND VPWR VGND VPWR _2734_ i_tinyqv.cpu.data_addr\[24\] _2853_ _1540_ sky130_fd_sc_hd__a21oi_2
Xi_tinyqv.cpu.i_core.i_instrret.i_regbuf\[5\] i_tinyqv.cpu.i_core.i_instrret.reg_buf\[5\]
+ i_tinyqv.cpu.i_core.i_instrret.register\[9\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_1_Right_1 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7398_ VPWR VGND _3651_ _3645_ i_tinyqv.cpu.instr_data_start\[8\] VPWR VGND sky130_fd_sc_hd__and2_1
X_6349_ VPWR VGND VGND VPWR _2790_ _1711_ _2789_ sky130_fd_sc_hd__or2_1
X_8019_ i_uart_rx.fsm_state\[2\] clknet_leaf_30_clk _0154_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_51_clk VGND VPWR clknet_3_1__leaf_clk clknet_leaf_51_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_0_19_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_27_12 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_3981_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.cmp _0744_ _0824_ _0833_ sky130_fd_sc_hd__o21a_1
X_5720_ VGND VPWR VGND VPWR i_debug_uart_tx.fsm_state\[0\] i_debug_uart_tx.fsm_state\[2\]
+ _2367_ _2368_ sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_42_clk VGND VPWR clknet_3_5__leaf_clk clknet_leaf_42_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_5651_ VGND VPWR VPWR VGND _2319_ _2318_ _2309_ i_tinyqv.cpu.instr_data\[3\]\[9\]
+ sky130_fd_sc_hd__mux2_1
X_5582_ VGND VPWR VGND VPWR _0146_ net160 _2263_ _2269_ _2240_ sky130_fd_sc_hd__o211a_1
X_8370_ i_tinyqv.cpu.data_read_n\[0\] clknet_leaf_21_clk _0469_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_2
X_4602_ VGND VPWR _1437_ _1431_ _1438_ _1436_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_4533_ VGND VPWR VPWR VGND _1372_ i_tinyqv.cpu.instr_data_in\[6\] _0838_ i_tinyqv.cpu.instr_data_in\[2\]
+ sky130_fd_sc_hd__mux2_1
X_7321_ VGND VPWR VPWR VGND _3590_ _3556_ _3454_ _2155_ _3384_ _3290_ sky130_fd_sc_hd__a32o_1
X_7252_ VPWR VGND VGND VPWR _3335_ _3532_ _3533_ sky130_fd_sc_hd__nor2_1
X_4464_ VGND VPWR VPWR VGND _1305_ debug_rd_r\[0\] debug_register_data i_spi.spi_dc
+ sky130_fd_sc_hd__mux2_1
X_6203_ VPWR VGND VPWR VGND i_tinyqv.cpu.i_core.mem_op\[2\] _2685_ _0878_ i_tinyqv.cpu.i_core.mem_op\[1\]
+ _2686_ sky130_fd_sc_hd__or4_1
X_4395_ VGND VPWR VPWR VGND _1238_ i_tinyqv.mem.qspi_data_buf\[9\] _1017_ i_tinyqv.cpu.instr_data_in\[9\]
+ sky130_fd_sc_hd__mux2_1
X_7183_ VGND VPWR VGND VPWR _3482_ _3331_ _3471_ _1491_ _3481_ sky130_fd_sc_hd__a211o_1
X_6134_ VPWR VGND VGND VPWR _2642_ _0653_ i_tinyqv.cpu.is_alu_imm sky130_fd_sc_hd__nand2_2
X_6065_ VGND VPWR _0297_ _2600_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5016_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[3\] _1779_ _1250_ sky130_fd_sc_hd__nand2_1
X_6967_ VPWR VGND _3290_ _3289_ VPWR VGND sky130_fd_sc_hd__buf_2
X_5918_ VGND VPWR _0240_ _2510_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6898_ VGND VPWR _0474_ _3256_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_33_clk VGND VPWR clknet_3_7__leaf_clk clknet_leaf_33_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_0_8_440 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5849_ VGND VPWR _2467_ _2468_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_8568_ VGND VPWR net1 uio_oe[3] VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_7519_ VPWR VGND VGND VPWR _2067_ _2073_ _0602_ sky130_fd_sc_hd__nor2_1
X_8499_ i_tinyqv.cpu.i_core.i_instrret.data\[1\] clknet_leaf_45_clk i_tinyqv.cpu.i_core.i_instrret.reg_buf\[5\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.i_regbuf\[11\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[11\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[15\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_24_clk VGND VPWR clknet_3_6__leaf_clk clknet_leaf_24_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_4180_ VGND VPWR i_tinyqv.cpu.alu_op\[2\] _1027_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_7870_ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[25\] clknet_leaf_53_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[25\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6821_ VGND VPWR VGND VPWR _0459_ _0784_ _3123_ _3194_ _3093_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_15_clk VGND VPWR clknet_3_2__leaf_clk clknet_leaf_15_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_6752_ VPWR VGND VPWR VGND _3124_ _3039_ _3132_ _2306_ _0906_ _3131_ sky130_fd_sc_hd__a221o_1
X_3964_ VGND VPWR VPWR VGND _0658_ _0816_ _0815_ sky130_fd_sc_hd__xor2_1
X_5703_ VPWR VGND VGND VPWR i_debug_uart_tx.cycle_counter\[0\] _2356_ _0989_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_633 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_6683_ VGND VPWR VGND VPWR _3069_ _3040_ _3067_ _3068_ _3047_ sky130_fd_sc_hd__o211a_1
X_3895_ VPWR VGND VPWR VGND _0745_ _0743_ _0746_ _0747_ sky130_fd_sc_hd__a21o_1
X_5634_ VPWR VGND _2309_ _2308_ VPWR VGND sky130_fd_sc_hd__buf_4
X_8422_ i_tinyqv.cpu.i_core.imm_lo\[0\] clknet_leaf_23_clk _0520_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_8353_ i_tinyqv.cpu.instr_data_start\[11\] clknet_leaf_33_clk _0452_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_13_210 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5565_ VPWR VGND _2259_ _2256_ i_uart_rx.cycle_counter\[9\] VPWR VGND sky130_fd_sc_hd__and2_1
Xhold100 net129 i_tinyqv.cpu.data_out\[20\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7304_ VPWR VGND VPWR VGND _2126_ _3349_ _3289_ _3577_ _3576_ sky130_fd_sc_hd__or4b_1
Xhold133 net162 i_spi.clock_divider\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5496_ VGND VPWR _2209_ i_uart_tx.cycle_counter\[4\] i_uart_tx.cycle_counter\[5\]
+ _2206_ VPWR VGND sky130_fd_sc_hd__and3_1
Xhold111 net140 i_tinyqv.cpu.data_out\[17\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_8284_ i_tinyqv.mem.qspi_data_buf\[24\] clknet_leaf_14_clk _0383_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
Xhold122 net151 i_tinyqv.mem.q_ctrl.addr\[4\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 net173 i_tinyqv.cpu.data_addr\[15\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_254 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_4516_ VPWR VGND VPWR VGND i_tinyqv.cpu.i_core.mie\[18\] _0944_ _1355_ _1228_ net15
+ _1354_ sky130_fd_sc_hd__a221o_1
Xhold166 net195 _0196_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 VGND VPWR net206 i_uart_tx.cycle_counter\[1\] VPWR VGND sky130_fd_sc_hd__buf_1
Xhold155 net184 i_spi.end_txn_reg VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4447_ VGND VPWR VPWR VGND _1290_ _1151_ _1149_ _1146_ sky130_fd_sc_hd__mux2_1
X_7235_ VPWR VGND VGND VPWR _3521_ _3474_ net190 _3510_ _0546_ sky130_fd_sc_hd__o22a_1
Xhold188 net217 i_tinyqv.cpu.i_core.i_instrret.data\[2\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 net228 i_tinyqv.cpu.i_core.mepc\[12\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7166_ VGND VPWR VPWR VGND _3468_ _3466_ _3467_ _1510_ sky130_fd_sc_hd__mux2_1
X_4378_ VGND VPWR VPWR VGND _1221_ i_tinyqv.cpu.instr_data_in\[13\] _0838_ i_tinyqv.cpu.instr_data_in\[9\]
+ sky130_fd_sc_hd__mux2_1
X_6117_ VPWR VGND VGND VPWR _2056_ _2596_ _2629_ sky130_fd_sc_hd__nor2_1
X_7097_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.imm_lo\[3\] _3360_ _3406_ _0523_ sky130_fd_sc_hd__o21a_1
X_6048_ VGND VPWR VPWR VGND _2590_ i_tinyqv.cpu.instr_data\[1\]\[14\] _2462_ _1720_
+ sky130_fd_sc_hd__mux2_1
X_7999_ i_uart_rx.cycle_counter\[3\] clknet_leaf_30_clk _0134_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_67_482 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5350_ VPWR VGND VGND VPWR _0840_ _2087_ _2066_ sky130_fd_sc_hd__nor2_2
X_5281_ VPWR VGND _2033_ _2031_ i_tinyqv.cpu.i_core.multiplier.accum\[15\] VPWR VGND
+ sky130_fd_sc_hd__and2_1
XFILLER_0_23_596 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4301_ VPWR VGND VGND VPWR _1092_ _1148_ _1147_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_246 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_4232_ VPWR VGND VGND VPWR _1048_ _1079_ _1078_ sky130_fd_sc_hd__nand2_1
X_7020_ VGND VPWR _3336_ _3337_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_4_clk VGND VPWR clknet_3_0__leaf_clk clknet_leaf_4_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_4163_ VGND VPWR VGND VPWR _1010_ _0994_ _1006_ _1009_ _0945_ sky130_fd_sc_hd__o211a_1
X_4094_ VPWR VGND VPWR VGND i_tinyqv.cpu.i_core.i_instrret.data\[0\] _0929_ _0941_
+ _0931_ i_tinyqv.cpu.i_core.cycle_count\[0\] _0940_ sky130_fd_sc_hd__a221o_1
X_7922_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[13\] clknet_leaf_25_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[13\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7853_ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[8\] clknet_leaf_49_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[8\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4996_ VPWR VGND VGND VPWR _1758_ _1759_ _1760_ sky130_fd_sc_hd__nor2_1
X_6804_ VPWR VGND VGND VPWR _3166_ _3179_ _3178_ sky130_fd_sc_hd__nand2_1
X_7784_ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[3\] clknet_leaf_57_clk _0077_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6735_ VPWR VGND VGND VPWR _3114_ _3116_ _3115_ sky130_fd_sc_hd__nand2_1
X_3947_ VGND VPWR VPWR VGND _0799_ _0798_ _0654_ _0788_ sky130_fd_sc_hd__mux2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.i_regbuf\[25\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[25\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[29\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6666_ VPWR VGND VGND VPWR i_tinyqv.cpu.instr_data_start\[5\] i_tinyqv.cpu.i_core.imm_lo\[5\]
+ _3053_ sky130_fd_sc_hd__nor2_1
X_3878_ VPWR VGND VPWR VGND _0642_ i_tinyqv.cpu.i_core.i_registers.reg_access\[12\]\[0\]
+ net74 _0730_ i_tinyqv.cpu.i_core.i_registers.reg_access\[9\]\[0\] sky130_fd_sc_hd__a22o_1
XFILLER_0_45_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5617_ VGND VPWR _2294_ _2296_ i_uart_rx.fsm_state\[3\] VPWR VGND sky130_fd_sc_hd__xnor2_1
X_8405_ i_tinyqv.cpu.data_out\[30\] clknet_leaf_20_clk _0503_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_6597_ VGND VPWR _2306_ _2995_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_5548_ _2246_ _2247_ _2248_ net17 VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_8336_ i_tinyqv.cpu.instr_write_offset\[1\] clknet_leaf_21_clk _0435_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_8267_ i_tinyqv.cpu.instr_data_in\[7\] clknet_leaf_14_clk _0366_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_2
X_5479_ VPWR VGND VPWR VGND _2197_ i_uart_tx.fsm_state\[0\] _0990_ sky130_fd_sc_hd__or2_2
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.i_regbuf\[14\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[14\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[18\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7218_ VPWR VGND _3511_ _3374_ _3330_ _3328_ _3362_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_8198_ i_tinyqv.cpu.i_core.i_shift.a\[17\] clknet_leaf_40_clk _0310_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_7149_ VPWR VGND VPWR VGND _3453_ _3452_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_493 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xclkbuf_3_7__f_clk VGND VPWR VGND VPWR clknet_0_clk clknet_3_7__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_4850_ VGND VPWR VPWR VGND _1666_ i_tinyqv.cpu.debug_rd\[1\] _1664_ i_tinyqv.cpu.i_core.i_registers.reg_access\[10\]\[1\]
+ sky130_fd_sc_hd__mux2_1
X_3801_ VPWR VGND _0653_ i_tinyqv.cpu.debug_instr_valid VPWR VGND sky130_fd_sc_hd__buf_4
X_6520_ VGND VPWR VPWR VGND _2933_ _2932_ _2920_ net11 sky130_fd_sc_hd__mux2_1
X_4781_ VPWR VGND VPWR VGND _0986_ i_spi.data\[7\] _1000_ _1616_ net9 sky130_fd_sc_hd__a22o_1
X_6451_ VPWR VGND VGND VPWR _2832_ _2880_ _2879_ sky130_fd_sc_hd__nand2_1
X_6382_ VGND VPWR VPWR VGND _2822_ _2821_ _2811_ i_tinyqv.mem.q_ctrl.read_cycles_count\[1\]
+ sky130_fd_sc_hd__mux2_1
X_5402_ VPWR VGND VGND VPWR _1426_ _2127_ _2132_ sky130_fd_sc_hd__nor2_1
X_8121_ i_spi.data\[4\] clknet_leaf_18_clk _0233_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5333_ VPWR VGND _2075_ _2074_ i_tinyqv.cpu.i_core.time_hi\[0\] VPWR VGND sky130_fd_sc_hd__and2_1
X_8052_ i_debug_uart_tx.fsm_state\[1\] clknet_leaf_30_clk _0187_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_5264_ VPWR VGND VGND VPWR _2015_ _2017_ _2016_ sky130_fd_sc_hd__nand2_1
X_5195_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[9\] _1950_ _1813_ sky130_fd_sc_hd__nand2_1
X_4215_ VGND VPWR VPWR VGND _1062_ i_tinyqv.cpu.i_core.i_shift.a\[17\] _1027_ i_tinyqv.cpu.i_core.i_shift.a\[14\]
+ sky130_fd_sc_hd__mux2_1
X_7003_ VGND VPWR VGND VPWR _3323_ _3287_ _3322_ _3284_ _3290_ sky130_fd_sc_hd__a211o_1
X_4146_ VPWR VGND _0993_ _0989_ _0969_ i_tinyqv.cpu.data_addr\[2\] _0992_ VGND VPWR
+ sky130_fd_sc_hd__a31o_1
X_4077_ VPWR VGND VGND VPWR _0924_ i_tinyqv.cpu.i_core.imm_lo\[8\] i_tinyqv.cpu.i_core.imm_lo\[9\]
+ sky130_fd_sc_hd__or2_1
X_7905_ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[28\] clknet_leaf_48_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[28\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7836_ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[23\] clknet_leaf_1_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[23\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.i_regbuf\[26\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[26\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[30\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4979_ VGND VPWR _1747_ gpio_out_sel\[4\] _1737_ _1742_ VPWR VGND sky130_fd_sc_hd__and3_1
X_7767_ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[18\] clknet_leaf_54_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[18\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6718_ VGND VPWR VPWR VGND _3101_ _3100_ _2993_ _3094_ sky130_fd_sc_hd__mux2_1
X_7698_ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[13\] clknet_leaf_56_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[13\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6649_ VPWR VGND _3037_ _3026_ VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_0_33_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.i_regbuf\[15\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[15\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[19\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_8319_ i_tinyqv.mem.q_ctrl.spi_in_buffer\[7\] clknet_leaf_16_clk _0418_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.i_regbuf\[14\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[14\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[18\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_cycles.i_regbuf\[12\] i_tinyqv.cpu.i_core.i_cycles.reg_buf\[12\]
+ i_tinyqv.cpu.i_core.i_cycles.register\[16\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4000_ VGND VPWR _0851_ i_tinyqv.cpu.is_load i_tinyqv.cpu.debug_instr_valid i_tinyqv.cpu.no_write_in_progress
+ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_46_77 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5951_ VGND VPWR VPWR VGND _2533_ _2532_ _2524_ net111 sky130_fd_sc_hd__mux2_1
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_4902_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_registers.rd\[2\] i_tinyqv.cpu.i_core.i_registers.rd\[3\]
+ _1695_ sky130_fd_sc_hd__nor2_1
X_5882_ VPWR VGND VGND VPWR net106 _2484_ i_tinyqv.cpu.instr_data_in\[1\] _2485_ _0229_
+ sky130_fd_sc_hd__o22a_1
X_4833_ VGND VPWR VPWR VGND _1656_ i_tinyqv.cpu.debug_rd\[2\] _1653_ net103 sky130_fd_sc_hd__mux2_1
X_7621_ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[0\] clknet_leaf_1_clk _0042_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_452 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_7552_ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[27\] clknet_leaf_46_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[27\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_614 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4764_ VGND VPWR VPWR VGND i_tinyqv.cpu.instr_data_start\[23\] _1599_ _1333_ sky130_fd_sc_hd__xor2_1
X_6503_ VGND VPWR VPWR VGND _2917_ _2915_ _2916_ net10 sky130_fd_sc_hd__mux2_1
X_7483_ VPWR VGND VGND VPWR i_tinyqv.cpu.data_addr\[21\] _2682_ _3722_ _3723_ sky130_fd_sc_hd__o21a_1
X_6434_ VGND VPWR VGND VPWR _0400_ _1707_ _2863_ _2866_ _2832_ sky130_fd_sc_hd__o211a_1
X_4695_ VPWR VGND _1531_ i_tinyqv.mem.qspi_data_byte_idx\[0\] _0864_ VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_31_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_6365_ VPWR VGND VGND VPWR _2806_ _2786_ _2784_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_6296_ VGND VPWR _0371_ _2757_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5316_ VPWR VGND VPWR VGND _2062_ _2057_ sky130_fd_sc_hd__inv_2
X_8104_ i_tinyqv.cpu.instr_data\[0\]\[4\] clknet_leaf_10_clk _0216_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_8035_ i_tinyqv.cpu.instr_data\[3\]\[13\] clknet_leaf_12_clk _0170_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5247_ VGND VPWR _1999_ _2000_ _1998_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_5178_ VPWR VGND _1934_ _1933_ _1932_ VPWR VGND sky130_fd_sc_hd__and2_1
X_4129_ VGND VPWR VPWR VGND _0976_ i_tinyqv.cpu.instr_data_in\[12\] _0838_ i_tinyqv.cpu.instr_data_in\[8\]
+ sky130_fd_sc_hd__mux2_1
X_7819_ i_tinyqv.cpu.i_core.i_registers.reg_access\[6\]\[2\] clknet_leaf_5_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[6\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_474 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_34_477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_15_691 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.i_regbuf\[30\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[30\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[2\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_16_58 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.i_regbuf\[26\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[26\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[30\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_13 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_80_561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_4480_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[1\] _1319_ _1250_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_447 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_6150_ VGND VPWR VPWR VGND _2655_ _2654_ _2645_ i_tinyqv.cpu.i_core.i_shift.b\[3\]
+ sky130_fd_sc_hd__mux2_1
X_5101_ VGND VPWR _1835_ _1832_ _1860_ _1834_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_6081_ VGND VPWR _0305_ _2608_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5032_ _1794_ _1769_ _1770_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_6983_ VGND VPWR _1455_ _3305_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_5934_ VGND VPWR VPWR VGND _2521_ i_tinyqv.cpu.i_core.mepc\[9\] _2106_ i_tinyqv.cpu.i_core.i_shift.a\[13\]
+ sky130_fd_sc_hd__mux2_1
X_5865_ VGND VPWR VPWR VGND _2477_ i_tinyqv.cpu.instr_data\[0\]\[9\] _2469_ _2318_
+ sky130_fd_sc_hd__mux2_1
X_4816_ VGND VPWR VPWR VGND _1646_ net32 _1642_ i_tinyqv.cpu.i_core.i_registers.reg_access\[14\]\[3\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_7604_ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[15\] clknet_leaf_1_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[15\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5796_ VPWR VGND VPWR VGND _1725_ _1004_ net220 _2428_ sky130_fd_sc_hd__a21o_1
X_7535_ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[10\] clknet_leaf_45_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[10\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4747_ VGND VPWR _1319_ _1581_ _1582_ _1318_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_7466_ VPWR VGND VPWR VGND _3697_ _0784_ i_tinyqv.cpu.instr_data_start\[19\] _3708_
+ sky130_fd_sc_hd__a21oi_1
X_4678_ VGND VPWR VPWR VGND _1514_ _1432_ _1513_ _1512_ sky130_fd_sc_hd__mux2_4
X_6417_ VPWR VGND VGND VPWR _1715_ _2803_ _2848_ _2851_ _2852_ sky130_fd_sc_hd__o22ai_1
X_7397_ VPWR VGND VGND VPWR _3650_ i_tinyqv.cpu.instr_data_start\[8\] _3645_ sky130_fd_sc_hd__or2_1
X_6348_ VGND VPWR _2789_ i_tinyqv.mem.q_ctrl.fsm_state\[1\] i_tinyqv.mem.q_ctrl.fsm_state\[2\]
+ _1707_ VPWR VGND sky130_fd_sc_hd__and3_1
X_6279_ VGND VPWR VPWR VGND _2749_ i_tinyqv.cpu.instr_data_in\[4\] _2744_ _1712_ sky130_fd_sc_hd__mux2_1
X_8018_ i_uart_rx.fsm_state\[1\] clknet_leaf_28_clk _0153_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.i_regbuf\[4\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[4\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[8\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_35 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_3980_ VGND VPWR VGND VPWR _0832_ _0827_ _0828_ _0830_ _0831_ sky130_fd_sc_hd__o211a_1
X_5650_ VGND VPWR i_tinyqv.cpu.instr_data_in\[9\] _2318_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xclkbuf_0_clk VGND VPWR VGND VPWR clk clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_4601_ VPWR VGND VPWR VGND _1437_ i_tinyqv.cpu.was_early_branch sky130_fd_sc_hd__inv_2
X_5581_ VPWR VGND VGND VPWR _2269_ i_uart_rx.recieved_data\[4\] _2264_ sky130_fd_sc_hd__or2_1
X_4532_ VGND VPWR VPWR VGND _1371_ i_tinyqv.mem.qspi_data_buf\[10\] _1017_ i_tinyqv.cpu.instr_data_in\[10\]
+ sky130_fd_sc_hd__mux2_1
X_7320_ VGND VPWR _0563_ _3589_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4463_ VGND VPWR _0051_ _1304_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7251_ VPWR VGND _3532_ _3427_ _3325_ VPWR VGND sky130_fd_sc_hd__and2_1
X_6202_ VPWR VGND VPWR VGND _0725_ i_tinyqv.cpu.i_core.mem_op\[0\] _2684_ _2685_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_68_64 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4394_ VGND VPWR VPWR VGND _1237_ _1236_ _1012_ _1221_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_15_Right_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7182_ VPWR VGND VGND VPWR _3481_ _3290_ _3455_ sky130_fd_sc_hd__or2_1
X_6133_ VPWR VGND VPWR VGND _2641_ _2640_ sky130_fd_sc_hd__inv_2
X_6064_ VGND VPWR VPWR VGND _2600_ i_tinyqv.cpu.i_core.i_shift.a\[8\] _2593_ i_tinyqv.cpu.i_core.i_shift.a\[4\]
+ sky130_fd_sc_hd__mux2_1
X_5015_ VPWR VGND VGND VPWR _1776_ _1778_ _1777_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_24_Right_24 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6966_ VPWR VGND VGND VPWR _1426_ _3289_ _1420_ sky130_fd_sc_hd__nor2_2
X_5917_ VGND VPWR VPWR VGND _2510_ _2509_ _2502_ i_tinyqv.cpu.data_addr\[3\] sky130_fd_sc_hd__mux2_1
X_6897_ VGND VPWR VPWR VGND _3256_ _2647_ _3254_ i_debug_uart_tx.uart_tx_data\[1\]
+ sky130_fd_sc_hd__mux2_1
X_5848_ VPWR VGND VPWR VGND _1406_ _2460_ i_tinyqv.cpu.instr_write_offset\[2\] _2467_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_36_539 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_8567_ VGND VPWR uio_oe[5] uio_oe[2] VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_5779_ VPWR VGND _0196_ _2414_ _2221_ net194 _2416_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_7518_ VGND VPWR _0601_ _3749_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8498_ i_tinyqv.cpu.i_core.i_instrret.data\[0\] clknet_leaf_39_clk i_tinyqv.cpu.i_core.i_instrret.reg_buf\[4\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7449_ VGND VPWR VPWR VGND _3694_ _3693_ _2681_ i_tinyqv.cpu.data_addr\[16\] sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_33_Right_33 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_10_Left_91 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_42_Right_42 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_79_480 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_13_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.i_regbuf\[29\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[29\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[1\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_51_Right_51 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_35_561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_35_583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_22_299 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_60_Right_60 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6820_ VPWR VGND VGND VPWR _3026_ _3194_ _3193_ sky130_fd_sc_hd__nand2_1
X_6751_ VGND VPWR VGND VPWR _3131_ _3040_ _3129_ _3130_ _3047_ sky130_fd_sc_hd__o211a_1
X_3963_ VGND VPWR VPWR VGND _0815_ _0814_ _0698_ net16 sky130_fd_sc_hd__mux2_1
X_5702_ VGND VPWR VGND VPWR _0180_ i_debug_uart_tx.uart_tx_data\[7\] _2330_ _2355_
+ _2299_ sky130_fd_sc_hd__o211a_1
X_6682_ VPWR VGND VGND VPWR _1390_ _3068_ _2515_ sky130_fd_sc_hd__nand2_1
X_3894_ VGND VPWR _0746_ _0721_ _0742_ _0722_ VPWR VGND sky130_fd_sc_hd__and3_1
X_5633_ VGND VPWR VGND VPWR _2308_ _2307_ _1406_ i_tinyqv.cpu.instr_write_offset\[2\]
+ i_tinyqv.cpu.i_core.i_cycles.rstn sky130_fd_sc_hd__and4_4
X_8421_ i_tinyqv.cpu.is_system clknet_leaf_7_clk _0519_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5564_ VGND VPWR _0139_ _2258_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8352_ i_tinyqv.cpu.instr_data_start\[10\] clknet_leaf_25_clk _0451_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
Xhold101 net130 i_tinyqv.cpu.data_out\[14\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7303_ VPWR VGND VPWR VGND _2123_ _3321_ _1426_ _3576_ sky130_fd_sc_hd__or3_1
X_4515_ VPWR VGND VPWR VGND i_tinyqv.cpu.i_core.mepc\[2\] net19 _1354_ _1349_ i_tinyqv.cpu.i_core.mstatus_mte
+ _1353_ sky130_fd_sc_hd__a221o_1
Xhold134 net163 _0203_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5495_ VPWR VGND VPWR VGND _2206_ net174 _2208_ _0120_ sky130_fd_sc_hd__a21oi_1
X_8283_ i_tinyqv.mem.data_from_read\[23\] clknet_leaf_17_clk _0382_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
Xhold123 net152 i_tinyqv.cpu.i_core.i_registers.reg_access\[6\]\[3\] VPWR VGND VGND
+ VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 net141 i_tinyqv.cpu.alu_op\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 net174 i_uart_tx.cycle_counter\[4\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 net185 _0199_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4446_ VPWR VGND VGND VPWR _1048_ _1289_ _1288_ sky130_fd_sc_hd__nand2_1
Xhold167 net196 i_tinyqv.cpu.instr_len\[2\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7234_ VGND VPWR _3428_ _3359_ _3521_ _3315_ VPWR VGND sky130_fd_sc_hd__o21ai_1
Xhold178 net207 i_uart_rx.recieved_data\[4\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4377_ VGND VPWR VPWR VGND _1220_ i_tinyqv.mem.qspi_data_buf\[29\] _0974_ i_tinyqv.mem.qspi_data_buf\[25\]
+ sky130_fd_sc_hd__mux2_1
Xhold189 net218 i_tinyqv.cpu.i_core.time_hi\[1\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7165_ VPWR VGND VGND VPWR _3467_ _3334_ _3319_ sky130_fd_sc_hd__or2_1
X_6116_ VGND VPWR VGND VPWR _2626_ _0798_ _1124_ _2628_ _2627_ sky130_fd_sc_hd__a2bb2o_1
X_7096_ VPWR VGND VPWR VGND _3377_ _3405_ _3400_ _3362_ _3406_ sky130_fd_sc_hd__or4_1
X_6047_ VGND VPWR _0290_ _2589_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7998_ i_uart_rx.cycle_counter\[2\] clknet_leaf_31_clk _0133_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_6949_ VGND VPWR VPWR VGND _0504_ _3273_ _3269_ _1589_ _3277_ net110 sky130_fd_sc_hd__a32o_1
XFILLER_0_24_509 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_40_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5280_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.multiplier.accum\[15\] _2031_ _2032_
+ sky130_fd_sc_hd__nor2_1
X_4300_ VGND VPWR VPWR VGND _1147_ _1146_ _1088_ _1145_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_9 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4231_ VGND VPWR VPWR VGND _1078_ _1075_ _1077_ _1059_ sky130_fd_sc_hd__mux2_1
X_4162_ VGND VPWR VGND VPWR _1009_ net14 _1007_ gpio_out_sel\[4\] _1008_ sky130_fd_sc_hd__a211o_1
X_4093_ VPWR VGND VPWR VGND _0938_ _0934_ _0939_ _0940_ sky130_fd_sc_hd__a21oi_1
X_7921_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[12\] clknet_leaf_36_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[12\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7852_ i_tinyqv.cpu.i_core.i_registers.reg_access\[5\]\[3\] clknet_leaf_45_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[7\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4995_ VPWR VGND VGND VPWR i_tinyqv.cpu.is_load _1759_ _1442_ sky130_fd_sc_hd__nand2_1
X_6803_ VPWR VGND VGND VPWR _3167_ _3178_ _3165_ sky130_fd_sc_hd__nand2_1
X_7783_ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[2\] clknet_leaf_54_clk _0076_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_494 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_6734_ VPWR VGND VGND VPWR _3115_ i_tinyqv.cpu.instr_data_start\[11\] i_tinyqv.cpu.i_core.imm_lo\[11\]
+ sky130_fd_sc_hd__or2_1
XFILLER_0_14_80 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_3946_ VPWR VGND VGND VPWR _0798_ _0797_ _0793_ sky130_fd_sc_hd__nor2_4
X_8404_ i_tinyqv.cpu.data_out\[29\] clknet_leaf_20_clk _0502_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_6665_ VPWR VGND _3052_ i_tinyqv.cpu.i_core.imm_lo\[5\] i_tinyqv.cpu.instr_data_start\[5\]
+ VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_60_114 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_3877_ VGND VPWR VPWR VGND _0727_ _0728_ _0723_ _0729_ sky130_fd_sc_hd__or3_2
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.i_regbuf\[18\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[18\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[22\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5616_ VGND VPWR VGND VPWR _2295_ _2229_ _2280_ _2238_ _0154_ _2294_ sky130_fd_sc_hd__a2111oi_1
X_6596_ VPWR VGND VPWR VGND _2992_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[9\]
+ _2987_ _2994_ _2993_ sky130_fd_sc_hd__a22o_1
X_8335_ i_tinyqv.mem.q_ctrl.delay_cycles_cfg\[2\] clknet_leaf_16_clk _0434_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5547_ VPWR VGND _2247_ net224 i_uart_rx.cycle_counter\[1\] net91 i_uart_rx.cycle_counter\[3\]
+ VGND VPWR sky130_fd_sc_hd__a31o_1
X_5478_ VGND VPWR VGND VPWR _0115_ i_debug_uart_tx.uart_tx_data\[7\] _2169_ _2196_
+ _2182_ sky130_fd_sc_hd__o211a_1
X_8266_ i_tinyqv.cpu.instr_data_in\[6\] clknet_leaf_14_clk _0365_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_4429_ VPWR VGND VGND VPWR _1092_ _1272_ _1271_ sky130_fd_sc_hd__nand2_1
X_7217_ VPWR VGND _3510_ _3509_ VPWR VGND sky130_fd_sc_hd__buf_2
X_8197_ i_tinyqv.cpu.i_core.i_shift.a\[16\] clknet_leaf_41_clk _0309_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_7148_ VPWR VGND VGND VPWR _3290_ _3452_ _3451_ sky130_fd_sc_hd__nand2_1
X_7079_ VPWR VGND VGND VPWR _3367_ i_tinyqv.cpu.instr_data\[1\]\[6\] _3365_ i_tinyqv.cpu.instr_data\[0\]\[6\]
+ _3390_ _3389_ sky130_fd_sc_hd__o221a_2
XFILLER_0_20_523 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4780_ VGND VPWR VPWR VGND _1615_ i_tinyqv.cpu.instr_data_in\[7\] _1012_ i_tinyqv.cpu.instr_data_in\[15\]
+ sky130_fd_sc_hd__mux2_1
X_3800_ VPWR VGND VPWR VGND _0641_ _0651_ _0636_ _0652_ sky130_fd_sc_hd__or3_4
XFILLER_0_55_475 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_6450_ VPWR VGND _2879_ _2878_ i_tinyqv.cpu.data_addr\[23\] i_tinyqv.cpu.data_addr\[24\]
+ _2855_ VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_42_136 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6381_ VPWR VGND VGND VPWR _2815_ _2819_ _2813_ _2820_ _2821_ sky130_fd_sc_hd__o22a_1
X_5401_ VPWR VGND VGND VPWR _1477_ _1488_ _2131_ sky130_fd_sc_hd__nor2_1
X_8120_ i_spi.data\[3\] clknet_leaf_18_clk _0232_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_233 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5332_ VPWR VGND VGND VPWR _1604_ _2073_ _2074_ sky130_fd_sc_hd__nor2_1
X_8051_ i_debug_uart_tx.fsm_state\[0\] clknet_leaf_30_clk _0186_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_2
X_5263_ VGND VPWR _1990_ _1987_ _2016_ _1989_ VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_75 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5194_ VGND VPWR VPWR VGND _1947_ _0025_ _1949_ sky130_fd_sc_hd__xor2_1
X_4214_ VGND VPWR VPWR VGND _1061_ i_tinyqv.cpu.i_core.i_shift.a\[16\] _1028_ _1060_
+ sky130_fd_sc_hd__mux2_1
X_7002_ VPWR VGND VGND VPWR _3321_ _3322_ _2118_ sky130_fd_sc_hd__nor2_2
X_4145_ VPWR VGND VGND VPWR _0985_ _0991_ _0992_ sky130_fd_sc_hd__nor2_1
X_4076_ VPWR VGND VPWR VGND i_tinyqv.cpu.i_core.imm_lo\[5\] i_tinyqv.cpu.i_core.imm_lo\[4\]
+ i_tinyqv.cpu.i_core.imm_lo\[7\] _0923_ sky130_fd_sc_hd__or3_1
X_7904_ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[27\] clknet_leaf_53_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[27\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7835_ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[22\] clknet_leaf_3_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[22\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_601 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_4978_ VPWR VGND VPWR VGND _1741_ net197 _1746_ _0011_ sky130_fd_sc_hd__a21o_1
X_7766_ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[17\] clknet_leaf_54_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[17\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.i_regbuf\[19\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[19\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[23\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6717_ VGND VPWR VPWR VGND _3100_ _3099_ _2990_ _2521_ sky130_fd_sc_hd__mux2_1
X_7697_ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[12\] clknet_leaf_2_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[12\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_3929_ VPWR VGND VGND VPWR _0763_ _0781_ _0780_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_626 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_6648_ VGND VPWR VGND VPWR _0444_ _0884_ _3027_ _3036_ _2061_ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_8318_ i_tinyqv.mem.q_ctrl.spi_in_buffer\[6\] clknet_leaf_16_clk _0417_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6579_ VGND VPWR _0430_ _2981_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8249_ i_tinyqv.mem.instr_active clknet_leaf_20_clk _0349_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.i_regbuf\[22\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[22\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[26\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_501 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.i_regbuf\[11\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[11\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[15\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_37_464 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_12_309 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_instrret.i_regbuf\[21\] i_tinyqv.cpu.i_core.i_instrret.reg_buf\[21\]
+ i_tinyqv.cpu.i_core.i_instrret.register\[25\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5950_ VGND VPWR VPWR VGND _2532_ i_tinyqv.cpu.i_core.mepc\[14\] _2107_ i_tinyqv.cpu.i_core.i_shift.a\[18\]
+ sky130_fd_sc_hd__mux2_1
X_4901_ VGND VPWR _0065_ _1694_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5881_ VPWR VGND VGND VPWR net100 _2484_ i_tinyqv.cpu.instr_data_in\[0\] _2485_ _0228_
+ sky130_fd_sc_hd__o22a_1
X_7620_ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[31\] clknet_leaf_2_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[31\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4832_ VGND VPWR _0039_ _1655_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4763_ VPWR VGND VPWR VGND _1594_ _1598_ _0688_ _1589_ _1590_ _1597_ sky130_fd_sc_hd__a2111o_1
X_7551_ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[26\] clknet_leaf_46_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[26\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6502_ VPWR VGND VGND VPWR _2916_ _2787_ _2795_ sky130_fd_sc_hd__nand2_2
X_4694_ VGND VPWR VGND VPWR _1530_ _1525_ _1521_ _0749_ _1529_ sky130_fd_sc_hd__o211ai_2
X_7482_ VPWR VGND VPWR VGND _3632_ _3219_ _3722_ _3719_ _3721_ _2877_ sky130_fd_sc_hd__a221o_1
XFILLER_0_16_648 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_6433_ VGND VPWR _2865_ _2863_ _2866_ _2853_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_6364_ VPWR VGND VGND VPWR _2787_ _2805_ _2799_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_6295_ VGND VPWR VPWR VGND _2757_ _1712_ _1552_ net293 sky130_fd_sc_hd__mux2_1
X_8103_ i_tinyqv.cpu.instr_data\[0\]\[3\] clknet_leaf_12_clk _0215_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5315_ _0087_ _2053_ _2058_ _2060_ _2061_ VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_0_53_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5246_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[12\] _1999_ _1880_ sky130_fd_sc_hd__nand2_1
X_8034_ i_tinyqv.cpu.instr_data\[3\]\[12\] clknet_leaf_11_clk _0169_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5177_ VPWR VGND VGND VPWR _1933_ _1928_ _1931_ sky130_fd_sc_hd__or2_1
X_4128_ VGND VPWR VPWR VGND _0975_ i_tinyqv.mem.qspi_data_buf\[28\] _0974_ i_tinyqv.mem.qspi_data_buf\[24\]
+ sky130_fd_sc_hd__mux2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.i_regbuf\[9\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[9\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[13\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4059_ VGND VPWR _0894_ _0906_ _0726_ VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_504 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_7818_ i_tinyqv.cpu.i_core.i_registers.reg_access\[6\]\[1\] clknet_leaf_5_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[5\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7749_ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[0\] clknet_leaf_57_clk _0078_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_191 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_30_640 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.i_regbuf\[23\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[23\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[27\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_16_37 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.i_regbuf\[19\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[19\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[23\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.i_regbuf\[12\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[12\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[16\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_228 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_80_551 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_52_231 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_501 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_5100_ VPWR VGND _1859_ _1858_ _1857_ VPWR VGND sky130_fd_sc_hd__and2_1
X_6080_ VGND VPWR VPWR VGND _2608_ i_tinyqv.cpu.i_core.i_shift.a\[16\] _2592_ i_tinyqv.cpu.i_core.i_shift.a\[12\]
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_29_Left_110 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5031_ VGND VPWR VPWR VGND _1791_ _1793_ _1792_ sky130_fd_sc_hd__xor2_1
X_6982_ VGND VPWR _1452_ _3304_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_5933_ VGND VPWR _0245_ _2520_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5864_ VGND VPWR _0220_ _2476_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_645 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_4815_ VGND VPWR _0048_ _1645_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7603_ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[14\] clknet_leaf_2_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[14\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5795_ VPWR VGND VGND VPWR _1004_ _2427_ _1725_ sky130_fd_sc_hd__nand2_1
X_7534_ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[9\] clknet_leaf_47_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[9\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4746_ VPWR VGND VGND VPWR _1581_ _1308_ _1317_ sky130_fd_sc_hd__or2_1
X_7465_ VGND VPWR _3707_ _0784_ i_tinyqv.cpu.instr_data_start\[19\] _3697_ VPWR VGND
+ sky130_fd_sc_hd__and3_1
X_4677_ VGND VPWR VPWR VGND _1513_ i_tinyqv.cpu.instr_data\[2\]\[8\] _1504_ i_tinyqv.cpu.instr_data\[0\]\[8\]
+ sky130_fd_sc_hd__mux2_1
X_6416_ VPWR VGND VPWR VGND _2851_ i_tinyqv.mem.q_ctrl.nibbles_remaining\[2\] sky130_fd_sc_hd__inv_2
X_7396_ VPWR VGND VGND VPWR _3625_ net302 _3624_ net95 _0579_ _3649_ sky130_fd_sc_hd__o221a_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.i_regbuf\[5\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[5\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[9\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6347_ VPWR VGND VGND VPWR _1713_ _2787_ _2788_ sky130_fd_sc_hd__nor2_1
X_6278_ VGND VPWR _0362_ _2748_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8017_ i_uart_rx.fsm_state\[0\] clknet_leaf_27_clk _0152_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_5229_ VPWR VGND _1983_ _1982_ _1981_ VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_22_415 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.i_regbuf\[4\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[4\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[8\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4600_ VPWR VGND _1436_ _1427_ _1432_ _1406_ _1435_ VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_26_710 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5580_ VGND VPWR VGND VPWR _0145_ net207 _2263_ _2268_ _2240_ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_359 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_25_220 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4531_ VGND VPWR VPWR VGND _1370_ i_tinyqv.mem.qspi_data_buf\[14\] _1017_ i_tinyqv.cpu.instr_data_in\[14\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_136 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_13_415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4462_ VGND VPWR VPWR VGND _1304_ i_tinyqv.cpu.debug_rd\[1\] _1190_ i_tinyqv.cpu.i_core.i_registers.reg_access\[15\]\[1\]
+ sky130_fd_sc_hd__mux2_1
X_7250_ VGND VPWR VGND VPWR _3531_ _3304_ _3315_ _3530_ _1493_ sky130_fd_sc_hd__o211a_1
X_6201_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.mem_op\[0\] _0939_ _2684_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_4393_ VGND VPWR VPWR VGND _1236_ i_tinyqv.cpu.instr_data_in\[5\] _0838_ i_tinyqv.cpu.instr_data_in\[1\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_331 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7181_ VPWR VGND VPWR VGND _3476_ _2124_ _3479_ _3480_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_386 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_6132_ VPWR VGND _0714_ _2640_ net59 VPWR VGND sky130_fd_sc_hd__and2_2
X_6063_ VGND VPWR _0296_ _2599_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5014_ VPWR VGND VGND VPWR _1765_ _1766_ _1777_ _1775_ sky130_fd_sc_hd__nand3_1
X_6965_ VPWR VGND VPWR VGND _3288_ _3287_ sky130_fd_sc_hd__inv_2
X_5916_ VGND VPWR VPWR VGND _2509_ i_tinyqv.cpu.i_core.mepc\[3\] _2106_ _1054_ sky130_fd_sc_hd__mux2_1
X_6896_ VGND VPWR _0473_ _3255_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5847_ VGND VPWR _0213_ _2466_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8566_ VGND VPWR uio_oe[5] uio_oe[1] VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_5778_ VPWR VGND VPWR VGND _2416_ _2415_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_242 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_8497_ i_tinyqv.mem.q_ctrl.addr\[23\] clknet_leaf_29_clk _0595_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_2
X_4729_ _1564_ _0823_ _1178_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_7517_ VGND VPWR VPWR VGND _3749_ _2644_ _3748_ i_tinyqv.cpu.i_core.i_shift.b\[4\]
+ sky130_fd_sc_hd__mux2_1
X_7448_ VGND VPWR _3169_ _3692_ _3693_ _1437_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_7379_ VPWR VGND VGND VPWR _3010_ _3634_ _3635_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_54_78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6750_ VPWR VGND VGND VPWR _1390_ _3130_ _2528_ sky130_fd_sc_hd__nand2_1
X_5701_ VPWR VGND VPWR VGND _2336_ net278 _2341_ _2355_ sky130_fd_sc_hd__a21o_1
X_3962_ VGND VPWR _0813_ _0752_ _0814_ _0810_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_6681_ VGND VPWR _3066_ _3067_ _3065_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_3893_ VGND VPWR VPWR VGND _0745_ _0658_ _0744_ i_tinyqv.cpu.i_core.cy sky130_fd_sc_hd__mux2_1
X_5632_ _2307_ _1552_ i_tinyqv.cpu.instr_fetch_running i_tinyqv.mem.instr_active _2306_
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
XFILLER_0_26_540 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_8420_ i_tinyqv.cpu.is_jal clknet_leaf_7_clk _0518_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_5563_ _2256_ _2242_ _2258_ _2257_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_8351_ i_tinyqv.cpu.instr_data_start\[9\] clknet_leaf_25_clk _0450_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_79_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7302_ VGND VPWR _0559_ _3575_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4514_ VGND VPWR VGND VPWR _1353_ _0929_ _1350_ i_tinyqv.cpu.i_core.i_instrret.data\[2\]
+ _1352_ sky130_fd_sc_hd__a211o_1
Xhold113 net142 i_uart_rx.cycle_counter\[10\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 net164 i_uart_tx.fsm_state\[2\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5494_ VGND VPWR _2206_ _2200_ _2208_ i_uart_tx.cycle_counter\[4\] VPWR VGND sky130_fd_sc_hd__o21ai_1
Xhold102 net131 i_tinyqv.cpu.data_out\[11\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 net153 i_tinyqv.mem.q_ctrl.addr\[8\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_8282_ i_tinyqv.mem.data_from_read\[22\] clknet_leaf_13_clk _0381_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
Xhold168 VGND VPWR net197 i_debug_uart_tx.uart_tx_data\[3\] VPWR VGND sky130_fd_sc_hd__buf_1
Xhold157 net186 i_spi.end_txn VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 net175 i_tinyqv.cpu.data_out\[18\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7233_ VGND VPWR _0545_ _3520_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4445_ VGND VPWR VPWR VGND _1288_ _1287_ _1077_ _1284_ sky130_fd_sc_hd__mux2_1
Xhold179 net208 i_tinyqv.mem.q_ctrl.spi_ram_a_select VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4376_ VPWR VGND VPWR VGND i_tinyqv.mem.data_from_read\[17\] _0689_ _1219_ _0748_
+ i_tinyqv.mem.data_from_read\[21\] _0957_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_7164_ VPWR VGND _3466_ _3374_ _1466_ _2155_ _3465_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_6115_ VPWR VGND VPWR VGND _2625_ net16 _0845_ _2627_ sky130_fd_sc_hd__a21oi_1
X_7095_ VPWR VGND VPWR VGND _3404_ _3364_ _3403_ _3405_ _2165_ sky130_fd_sc_hd__a22o_1
X_6046_ VGND VPWR VPWR VGND _2589_ i_tinyqv.cpu.instr_data\[1\]\[13\] _2462_ _1717_
+ sky130_fd_sc_hd__mux2_1
X_7997_ i_uart_rx.cycle_counter\[1\] clknet_leaf_30_clk _0132_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_6948_ VGND VPWR VPWR VGND _0503_ _3273_ _3268_ _1589_ _3277_ net120 sky130_fd_sc_hd__a32o_1
X_6879_ VGND VPWR VGND VPWR _0467_ _1762_ _3244_ i_tinyqv.cpu.i_core.mem_op\[0\] _2067_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_48_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_551 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_8549_ i_tinyqv.cpu.i_core.i_cycles.register\[22\] clknet_leaf_4_clk i_tinyqv.cpu.i_core.i_cycles.reg_buf\[22\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_24_37 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4230_ VGND VPWR _1076_ _1077_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_4161_ VPWR VGND VPWR VGND _1001_ i_spi.data\[4\] _1000_ _1008_ uo_out[4] sky130_fd_sc_hd__a22o_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.i_regbuf\[26\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[26\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[30\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4092_ VPWR VGND VGND VPWR _0748_ _0939_ _0752_ sky130_fd_sc_hd__nand2_4
X_7920_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[11\] clknet_leaf_24_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[11\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7851_ i_tinyqv.cpu.i_core.i_registers.reg_access\[5\]\[2\] clknet_leaf_5_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[6\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6802_ VPWR VGND VGND VPWR _3175_ _3177_ _3176_ sky130_fd_sc_hd__nand2_1
X_7782_ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[1\] clknet_leaf_55_clk _0075_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4994_ VPWR VGND _1758_ _1757_ VPWR VGND sky130_fd_sc_hd__buf_4
XFILLER_0_46_602 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_6733_ VPWR VGND VGND VPWR i_tinyqv.cpu.instr_data_start\[11\] _3114_ i_tinyqv.cpu.i_core.imm_lo\[11\]
+ sky130_fd_sc_hd__nand2_1
X_3945_ VGND VPWR VGND VPWR _0649_ i_tinyqv.cpu.i_core.i_registers.reg_access\[7\]\[2\]
+ _0794_ _0795_ _0797_ _0796_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_45_101 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_6664_ VGND VPWR _2993_ _3051_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_5615_ VGND VPWR VGND VPWR i_uart_rx.fsm_state\[2\] _2289_ _2292_ _2295_ sky130_fd_sc_hd__o21ba_1
X_8403_ i_tinyqv.cpu.data_out\[28\] clknet_leaf_20_clk _0501_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_3876_ VGND VPWR VPWR VGND _0728_ _0619_ _0611_ i_tinyqv.cpu.instr_data_start\[4\]
+ _0613_ i_tinyqv.cpu.instr_data_start\[16\] sky130_fd_sc_hd__a32o_1
X_6595_ VGND VPWR net40 _2993_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_54_690 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_8334_ i_tinyqv.mem.q_ctrl.delay_cycles_cfg\[1\] clknet_leaf_15_clk _0433_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5546_ VGND VPWR _2246_ i_uart_rx.cycle_counter\[2\] i_uart_rx.cycle_counter\[3\]
+ _2236_ VPWR VGND sky130_fd_sc_hd__and3_1
X_5477_ VPWR VGND VPWR VGND _2195_ i_uart_tx.data_to_send\[7\] _2179_ _2196_ sky130_fd_sc_hd__a21o_1
X_8265_ i_tinyqv.cpu.instr_data_in\[5\] clknet_leaf_14_clk _0364_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_2
X_4428_ VGND VPWR VPWR VGND _1271_ _1070_ _1149_ _1066_ sky130_fd_sc_hd__mux2_1
X_7216_ VPWR VGND VPWR VGND _3464_ _3363_ _3499_ _3509_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_481 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_8196_ i_tinyqv.cpu.i_core.i_shift.a\[15\] clknet_leaf_41_clk _0308_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_4359_ VGND VPWR VPWR VGND _0882_ _1202_ _0892_ sky130_fd_sc_hd__xor2_1
X_7147_ VPWR VGND VGND VPWR _3368_ i_tinyqv.cpu.instr_data\[1\]\[13\] _3366_ i_tinyqv.cpu.instr_data\[0\]\[13\]
+ _3451_ _3450_ sky130_fd_sc_hd__o221a_1
X_7078_ VPWR VGND VPWR VGND i_tinyqv.cpu.instr_data\[3\]\[6\] _1504_ _3389_ _1461_
+ i_tinyqv.cpu.instr_data\[2\]\[6\] _3371_ sky130_fd_sc_hd__a221o_1
X_6029_ VGND VPWR _0281_ _2580_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xi_tinyqv.cpu.i_core.i_cycles.i_regbuf\[9\] i_tinyqv.cpu.i_core.i_cycles.reg_buf\[9\]
+ i_tinyqv.cpu.i_core.i_cycles.register\[13\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_395 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_20_579 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_27_178 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_6380_ VPWR VGND _2820_ _2784_ i_tinyqv.mem.q_ctrl.delay_cycles_cfg\[2\] _2792_ _2787_
+ VGND VPWR sky130_fd_sc_hd__a31o_1
X_5400_ VGND VPWR VGND VPWR _2129_ _2130_ _2122_ _2123_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_42_159 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_5331_ VPWR VGND VGND VPWR net235 _2073_ _2072_ sky130_fd_sc_hd__nand2_1
X_8050_ i_debug_uart_tx.cycle_counter\[4\] clknet_leaf_30_clk _0185_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.i_regbuf\[27\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[27\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[31\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5262_ VGND VPWR VPWR VGND _2013_ _2015_ _2014_ sky130_fd_sc_hd__xor2_1
X_7001_ VPWR VGND VGND VPWR _1420_ _3321_ _1476_ sky130_fd_sc_hd__nand2_1
X_5193_ VPWR VGND VGND VPWR _1919_ _1949_ _1948_ sky130_fd_sc_hd__nand2_1
X_4213_ VPWR VGND _1060_ i_tinyqv.cpu.i_core.i_shift.a\[15\] VPWR VGND sky130_fd_sc_hd__buf_2
X_4144_ VPWR VGND VGND VPWR _0991_ _0990_ i_uart_tx.fsm_state\[0\] sky130_fd_sc_hd__nor2_4
X_4075_ VPWR VGND VPWR VGND i_tinyqv.cpu.i_core.imm_lo\[1\] i_tinyqv.cpu.i_core.imm_lo\[0\]
+ _0922_ i_tinyqv.cpu.i_core.imm_lo\[3\] i_tinyqv.cpu.i_core.imm_lo\[2\] sky130_fd_sc_hd__or4b_2
X_7903_ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[26\] clknet_leaf_3_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[26\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7834_ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[21\] clknet_leaf_3_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[21\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.i_regbuf\[30\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[30\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[2\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7765_ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[16\] clknet_leaf_1_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[16\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_613 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4977_ VGND VPWR _1746_ gpio_out_sel\[3\] _1737_ _1742_ VPWR VGND sky130_fd_sc_hd__and3_1
X_6716_ VGND VPWR VPWR VGND _3095_ _3099_ _3098_ sky130_fd_sc_hd__xor2_1
XFILLER_0_73_262 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7696_ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[11\] clknet_leaf_57_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[11\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_679 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_3928_ VGND VPWR VPWR VGND _0658_ _0780_ _0779_ sky130_fd_sc_hd__xor2_1
X_6647_ VPWR VGND VGND VPWR _3036_ _3029_ _3035_ sky130_fd_sc_hd__or2_1
X_3859_ VPWR VGND _0711_ _0663_ _0662_ VPWR VGND sky130_fd_sc_hd__and2_1
X_6578_ VGND VPWR VPWR VGND _2981_ _2980_ _2562_ i_tinyqv.cpu.instr_data_in\[0\] sky130_fd_sc_hd__mux2_1
XFILLER_0_6_584 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_8317_ i_tinyqv.mem.q_ctrl.spi_in_buffer\[5\] clknet_leaf_16_clk _0416_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5529_ VGND VPWR i_uart_tx.fsm_state\[0\] _2233_ i_uart_tx.fsm_state\[2\] VPWR VGND
+ sky130_fd_sc_hd__xnor2_1
X_8248_ i_tinyqv.cpu.i_core.mepc\[19\] clknet_leaf_35_clk _0348_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_8179_ i_tinyqv.cpu.instr_data\[1\]\[14\] clknet_leaf_11_clk _0291_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.i_regbuf\[15\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[15\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[19\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_49_281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_24_159 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_33_682 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_20_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xi_tinyqv.cpu.i_core.i_instrret.i_regbuf\[14\] i_tinyqv.cpu.i_core.i_instrret.reg_buf\[14\]
+ i_tinyqv.cpu.i_core.i_instrret.register\[18\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_5880_ VPWR VGND _2485_ _2307_ _1406_ i_tinyqv.cpu.instr_write_offset\[2\] _2066_
+ VGND VPWR sky130_fd_sc_hd__a31o_1
X_4900_ VGND VPWR VPWR VGND _1694_ _1638_ _1690_ i_tinyqv.cpu.i_core.i_registers.reg_access\[5\]\[3\]
+ sky130_fd_sc_hd__mux2_1
X_4831_ VGND VPWR VPWR VGND _1655_ i_tinyqv.cpu.debug_rd\[1\] _1653_ i_tinyqv.cpu.i_core.i_registers.reg_access\[12\]\[1\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_4762_ VPWR VGND VGND VPWR _0909_ _1596_ _1597_ sky130_fd_sc_hd__nor2_1
X_7550_ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[25\] clknet_leaf_54_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[25\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6501_ VGND VPWR VPWR VGND _2915_ _2913_ _2914_ _2910_ sky130_fd_sc_hd__mux2_1
X_4693_ VPWR VGND VPWR VGND _1528_ _1529_ net60 _1524_ sky130_fd_sc_hd__a21boi_1
X_7481_ VPWR VGND VGND VPWR _3010_ _3720_ _3721_ sky130_fd_sc_hd__nor2_1
X_6432_ VGND VPWR VGND VPWR _2865_ _1707_ _2845_ _2864_ _2801_ sky130_fd_sc_hd__o211a_1
X_6363_ VPWR VGND VGND VPWR _2794_ _2803_ _2804_ sky130_fd_sc_hd__nor2_1
X_8102_ i_tinyqv.cpu.instr_data\[0\]\[2\] clknet_leaf_11_clk _0214_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_6294_ VGND VPWR _0370_ _2756_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5314_ VGND VPWR _1752_ _2061_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_8033_ i_tinyqv.cpu.instr_data\[3\]\[11\] clknet_leaf_11_clk _0168_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5245_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[11\] _1998_ _1813_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5176_ VPWR VGND VGND VPWR _1928_ _1932_ _1931_ sky130_fd_sc_hd__nand2_1
X_4127_ VPWR VGND _0974_ _0838_ VPWR VGND sky130_fd_sc_hd__buf_4
X_4058_ VPWR VGND VGND VPWR _0905_ _0889_ _0904_ sky130_fd_sc_hd__or2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.i_regbuf\[31\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[31\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[3\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_590 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_7817_ i_tinyqv.cpu.i_core.i_registers.reg_access\[6\]\[0\] clknet_leaf_49_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[4\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7748_ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[31\] clknet_leaf_55_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[31\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7679_ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[26\] clknet_leaf_58_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[26\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_402 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.i_regbuf\[20\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[20\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[24\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.i_regbuf\[27\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[27\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[31\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.i_regbuf\[16\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[16\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[20\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_54_clk VGND VPWR clknet_3_1__leaf_clk clknet_leaf_54_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_0_37_240 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_557 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5030_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[5\] _1792_ _1166_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_129 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6981_ VGND VPWR VGND VPWR _3303_ _2123_ _2122_ _3297_ _3302_ sky130_fd_sc_hd__o211a_1
X_5932_ VGND VPWR VPWR VGND _2520_ _2519_ _2502_ i_tinyqv.cpu.data_addr\[8\] sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_45_clk VGND VPWR clknet_3_4__leaf_clk clknet_leaf_45_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_0_48_516 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_5863_ VGND VPWR VPWR VGND _2476_ i_tinyqv.cpu.instr_data\[0\]\[8\] _2469_ _2316_
+ sky130_fd_sc_hd__mux2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.i_regbuf\[7\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[7\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[11\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5794_ VGND VPWR _0201_ _2426_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4814_ VGND VPWR VPWR VGND _1645_ i_tinyqv.cpu.debug_rd\[2\] _1642_ i_tinyqv.cpu.i_core.i_registers.reg_access\[14\]\[2\]
+ sky130_fd_sc_hd__mux2_1
X_7602_ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[13\] clknet_leaf_53_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[13\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_571 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_7533_ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[8\] clknet_leaf_46_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[8\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4745_ VGND VPWR VPWR VGND _1578_ _1580_ _1579_ sky130_fd_sc_hd__xor2_1
X_7464_ VPWR VGND VGND VPWR net189 _3625_ _3706_ _0590_ sky130_fd_sc_hd__o21a_1
XFILLER_0_43_287 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4676_ VGND VPWR VPWR VGND _1512_ i_tinyqv.cpu.instr_data\[3\]\[8\] _1504_ i_tinyqv.cpu.instr_data\[1\]\[8\]
+ sky130_fd_sc_hd__mux2_1
X_6415_ VGND VPWR VPWR VGND _0397_ _2844_ _2832_ net265 _2850_ _2811_ sky130_fd_sc_hd__a32o_1
X_7395_ VGND VPWR VGND VPWR _3649_ _2878_ _2733_ net297 _3648_ sky130_fd_sc_hd__a211o_1
X_6346_ VPWR VGND _2787_ _2786_ VPWR VGND sky130_fd_sc_hd__buf_2
X_8016_ i_uart_rx.uart_rts clknet_leaf_27_clk _0151_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6277_ VGND VPWR VPWR VGND _2748_ i_tinyqv.cpu.instr_data_in\[3\] _2744_ _2322_ sky130_fd_sc_hd__mux2_1
X_5228_ VPWR VGND VGND VPWR _1982_ _1978_ _1980_ sky130_fd_sc_hd__or2_1
X_5159_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[9\] _1916_ _1845_ sky130_fd_sc_hd__nand2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.i_regbuf\[5\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[5\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[9\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_36_clk VGND VPWR clknet_3_6__leaf_clk clknet_leaf_36_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.i_regbuf\[31\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[31\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[3\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_27_clk VGND VPWR clknet_3_6__leaf_clk clknet_leaf_27_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_4530_ VGND VPWR VGND VPWR _1369_ _1364_ _1365_ _1368_ _0945_ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_202 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4461_ VPWR VGND i_tinyqv.cpu.debug_rd\[1\] _1303_ VPWR VGND sky130_fd_sc_hd__buf_2
X_6200_ VPWR VGND _2683_ _1026_ i_tinyqv.cpu.i_core.load_top_bit VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_40_246 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_7180_ VPWR VGND VPWR VGND _3465_ _3315_ _2140_ _3479_ sky130_fd_sc_hd__a21o_1
X_4392_ VGND VPWR VPWR VGND _1235_ i_tinyqv.mem.qspi_data_buf\[13\] _1017_ i_tinyqv.cpu.instr_data_in\[13\]
+ sky130_fd_sc_hd__mux2_1
X_6131_ VGND VPWR _0324_ _2639_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_365 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6062_ VGND VPWR VPWR VGND _2599_ _1054_ _2593_ i_tinyqv.cpu.i_core.i_shift.a\[3\]
+ sky130_fd_sc_hd__mux2_1
X_5013_ VPWR VGND VPWR VGND _1766_ _1765_ _1775_ _1776_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_18_clk VGND VPWR clknet_3_3__leaf_clk clknet_leaf_18_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_6964_ VGND VPWR VPWR VGND _3287_ _1432_ _3286_ _3285_ sky130_fd_sc_hd__mux2_4
XPHY_EDGE_ROW_5_Right_5 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6895_ VGND VPWR VPWR VGND _3255_ _2641_ _3254_ i_debug_uart_tx.uart_tx_data\[0\]
+ sky130_fd_sc_hd__mux2_1
X_5915_ VGND VPWR _0239_ _2508_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5846_ VGND VPWR VPWR VGND _2466_ _2465_ _2463_ i_tinyqv.cpu.instr_data_in\[1\] sky130_fd_sc_hd__mux2_1
XFILLER_0_8_421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_8565_ VGND VPWR net1 uio_oe[0] VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_5777_ VPWR VGND VGND VPWR _2415_ _1728_ _2394_ sky130_fd_sc_hd__nand2_2
X_8496_ i_tinyqv.mem.q_ctrl.addr\[22\] clknet_leaf_32_clk _0594_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_31_202 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4728_ VPWR VGND VGND VPWR _1563_ _0656_ i_tinyqv.cpu.alu_op\[3\] sky130_fd_sc_hd__nand2_2
X_7516_ VPWR VGND VGND VPWR _0939_ _1755_ _3748_ sky130_fd_sc_hd__nor2_1
X_7447_ VPWR VGND VPWR VGND _3690_ _3691_ i_tinyqv.cpu.was_early_branch _3692_ sky130_fd_sc_hd__or3_1
X_4659_ VGND VPWR VGND VPWR _1494_ _1490_ _1495_ sky130_fd_sc_hd__or2_4
XFILLER_0_31_268 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7378_ VGND VPWR VGND VPWR _3634_ i_tinyqv.cpu.instr_write_offset\[3\] _0884_ i_tinyqv.cpu.instr_data_start\[4\]
+ i_tinyqv.cpu.instr_data_start\[5\] sky130_fd_sc_hd__and4_2
X_6329_ VGND VPWR VPWR VGND _2776_ _2322_ _2772_ net253 sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_48_Left_129 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_57_Left_138 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_38_25 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_66_Left_147 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_3961_ VPWR VGND VGND VPWR _0813_ _0811_ _0812_ sky130_fd_sc_hd__or2_1
X_5700_ VGND VPWR VGND VPWR _0179_ net319 _2330_ _2354_ _2299_ sky130_fd_sc_hd__o211a_1
X_6680_ VGND VPWR VGND VPWR _3052_ _3053_ _3055_ _3066_ sky130_fd_sc_hd__o21ba_1
X_3892_ VPWR VGND VGND VPWR _0744_ _0612_ _0688_ sky130_fd_sc_hd__nor2_4
XPHY_EDGE_ROW_75_Left_156 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5631_ VPWR VGND VGND VPWR _2306_ _1546_ _1399_ sky130_fd_sc_hd__nor2_4
X_5562_ VPWR VGND _2257_ _2251_ i_uart_rx.cycle_counter\[6\] i_uart_rx.cycle_counter\[7\]
+ i_uart_rx.cycle_counter\[8\] VGND VPWR sky130_fd_sc_hd__a31o_1
X_8350_ i_tinyqv.cpu.instr_data_start\[8\] clknet_leaf_33_clk _0449_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
X_8281_ i_tinyqv.mem.data_from_read\[21\] clknet_leaf_13_clk _0380_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_7301_ VGND VPWR VPWR VGND _3575_ _3574_ _3395_ _0627_ sky130_fd_sc_hd__mux2_1
X_4513_ VPWR VGND VPWR VGND _1351_ i_tinyqv.cpu.i_core.cycle_count\[2\] _0931_ _1352_
+ _0927_ sky130_fd_sc_hd__a22o_1
Xhold103 net132 i_tinyqv.cpu.data_out\[10\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5493_ VPWR VGND VGND VPWR _2206_ _2207_ _0119_ sky130_fd_sc_hd__nor2_1
Xhold114 net143 i_tinyqv.cpu.data_out\[19\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7232_ VGND VPWR VPWR VGND _3520_ _3519_ _3396_ i_tinyqv.cpu.imm\[25\] sky130_fd_sc_hd__mux2_1
Xhold125 net154 i_tinyqv.cpu.additional_mem_ops\[2\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 net165 _2232_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 net187 i_tinyqv.mem.q_ctrl.addr\[9\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold147 net176 i_tinyqv.cpu.i_core.i_instrret.data\[1\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4444_ VGND VPWR VPWR VGND _1287_ _1286_ _1058_ _1285_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_7_clk VGND VPWR clknet_3_3__leaf_clk clknet_leaf_7_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold169 net198 i_tinyqv.cpu.i_core.i_registers.reg_access\[1\]\[0\] VPWR VGND VGND
+ VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4375_ VPWR VGND VGND VPWR _0878_ _1218_ _1217_ sky130_fd_sc_hd__nand2_1
X_7163_ VPWR VGND _3465_ _3464_ _1467_ VPWR VGND sky130_fd_sc_hd__and2_1
X_6114_ VPWR VGND VGND VPWR _2626_ _1326_ _1328_ _2625_ sky130_fd_sc_hd__nand3b_1
X_7094_ VPWR VGND VPWR VGND _3337_ _3350_ _3292_ _3404_ sky130_fd_sc_hd__or3_1
X_6045_ VGND VPWR _0289_ _2588_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7996_ i_uart_rx.cycle_counter\[0\] clknet_leaf_31_clk _0131_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_611 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6947_ VGND VPWR VPWR VGND _0502_ _3274_ _3267_ _1589_ _3277_ net109 sky130_fd_sc_hd__a32o_1
X_6878_ VPWR VGND VGND VPWR i_tinyqv.cpu.data_write_n\[0\] _1556_ _3243_ _3244_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_240 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5829_ VPWR VGND VGND VPWR net182 _2454_ _2453_ sky130_fd_sc_hd__nand2_1
X_8548_ i_tinyqv.cpu.i_core.i_cycles.register\[21\] clknet_leaf_3_clk i_tinyqv.cpu.i_core.i_cycles.reg_buf\[21\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_8479_ i_tinyqv.mem.q_ctrl.addr\[5\] clknet_leaf_32_clk _0577_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_588 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xi_tinyqv.cpu.i_core.i_cycles.i_regbuf\[28\] i_tinyqv.cpu.i_core.i_cycles.reg_buf\[28\]
+ i_tinyqv.cpu.i_core.i_cycles.register\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4160_ VPWR VGND VPWR VGND net6 _0986_ _1007_ _0997_ i_uart_rx.recieved_data\[4\]
+ _0908_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.i_regbuf\[19\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[19\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[23\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4091_ VPWR VGND VPWR VGND _0928_ _0937_ _0935_ _0938_ sky130_fd_sc_hd__or3_1
X_7850_ i_tinyqv.cpu.i_core.i_registers.reg_access\[5\]\[1\] clknet_leaf_47_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[5\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6801_ VPWR VGND VGND VPWR _3176_ i_tinyqv.cpu.instr_data_start\[17\] i_tinyqv.cpu.imm\[17\]
+ sky130_fd_sc_hd__or2_1
XFILLER_0_58_441 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7781_ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[0\] clknet_leaf_56_clk _0074_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4993_ VPWR VGND VGND VPWR _1757_ _0836_ _1756_ sky130_fd_sc_hd__or2_1
X_6732_ VGND VPWR VPWR VGND _3113_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[19\]
+ net31 _1596_ sky130_fd_sc_hd__mux2_1
X_3944_ VPWR VGND VPWR VGND _0642_ i_tinyqv.cpu.i_core.i_registers.reg_access\[5\]\[2\]
+ _0645_ _0796_ i_tinyqv.cpu.i_core.i_registers.reg_access\[9\]\[2\] sky130_fd_sc_hd__a22o_1
XFILLER_0_46_614 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6663_ VGND VPWR VGND VPWR _0445_ i_tinyqv.cpu.instr_data_start\[4\] _3027_ _3050_
+ _2061_ sky130_fd_sc_hd__o211a_1
X_3875_ VPWR VGND VPWR VGND _0725_ i_tinyqv.cpu.instr_data_start\[20\] _0610_ _0727_
+ _0726_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5614_ VGND VPWR _2294_ i_uart_rx.fsm_state\[1\] i_uart_rx.fsm_state\[2\] i_uart_rx.fsm_state\[0\]
+ VPWR VGND sky130_fd_sc_hd__and3_1
X_8402_ i_tinyqv.cpu.data_out\[27\] clknet_leaf_26_clk _0500_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_6594_ VGND VPWR VPWR VGND _2992_ _2988_ _2991_ _2505_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_533 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_8333_ i_tinyqv.mem.q_ctrl.delay_cycles_cfg\[0\] clknet_leaf_18_clk _0432_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5545_ VPWR VGND VPWR VGND _2236_ net178 _2245_ _0133_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5476_ VPWR VGND VPWR VGND _2195_ _2177_ sky130_fd_sc_hd__inv_2
X_8264_ i_tinyqv.cpu.instr_data_in\[4\] clknet_leaf_14_clk _0363_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_7215_ VPWR VGND VGND VPWR _3508_ _3474_ i_tinyqv.cpu.imm\[19\] _3500_ _0539_ sky130_fd_sc_hd__o22a_1
X_4427_ VGND VPWR VGND VPWR _1048_ _1269_ _1077_ _1263_ _1265_ _1270_ sky130_fd_sc_hd__a311o_1
X_8195_ i_tinyqv.cpu.i_core.i_shift.a\[14\] clknet_leaf_40_clk _0307_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
X_7146_ VPWR VGND VPWR VGND i_tinyqv.cpu.instr_data\[3\]\[13\] _3369_ _3450_ _3370_
+ i_tinyqv.cpu.instr_data\[2\]\[13\] _3372_ sky130_fd_sc_hd__a221o_1
X_4358_ VPWR VGND VGND VPWR _1201_ _0895_ _1200_ sky130_fd_sc_hd__or2_1
X_4289_ VGND VPWR VPWR VGND _1136_ _1135_ _1108_ _1134_ sky130_fd_sc_hd__mux2_1
X_7077_ VPWR VGND VGND VPWR _1491_ _3377_ _3348_ _3388_ sky130_fd_sc_hd__o21a_1
X_6028_ VGND VPWR VPWR VGND _2580_ i_tinyqv.cpu.instr_data\[1\]\[4\] _2463_ i_tinyqv.cpu.instr_data_in\[4\]
+ sky130_fd_sc_hd__mux2_1
X_7979_ i_uart_tx.data_to_send\[6\] clknet_leaf_28_clk _0114_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_488 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_44_190 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_60_661 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_19_49 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5330_ VGND VPWR _2072_ i_tinyqv.cpu.i_core.cycle_count\[1\] i_tinyqv.cpu.i_core.cycle_count\[2\]
+ _2071_ VPWR VGND sky130_fd_sc_hd__and3_1
X_5261_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[13\] _2014_ _1845_ sky130_fd_sc_hd__nand2_1
X_4212_ VGND VPWR VPWR VGND _1059_ _1056_ _1058_ _1052_ sky130_fd_sc_hd__mux2_1
X_7000_ VPWR VGND VGND VPWR _3305_ _3319_ _3320_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_44 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5192_ VGND VPWR VGND VPWR _1948_ _1922_ _1897_ _1921_ sky130_fd_sc_hd__a21bo_1
X_4143_ VPWR VGND VPWR VGND i_uart_tx.fsm_state\[2\] i_uart_tx.fsm_state\[1\] i_uart_tx.fsm_state\[3\]
+ _0990_ sky130_fd_sc_hd__or3_4
X_4074_ VPWR VGND _0921_ _0920_ _0858_ VPWR VGND sky130_fd_sc_hd__and2_1
X_7902_ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[25\] clknet_leaf_2_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[25\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7833_ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[20\] clknet_leaf_48_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[20\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7764_ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[15\] clknet_leaf_58_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[15\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4976_ VPWR VGND VPWR VGND _1741_ net98 _1745_ _0010_ sky130_fd_sc_hd__a21o_1
X_6715_ VPWR VGND VGND VPWR _3096_ _3098_ _3097_ sky130_fd_sc_hd__nand2_1
X_7695_ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[10\] clknet_leaf_53_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[10\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.i_regbuf\[23\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[23\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[27\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3927_ VPWR VGND VGND VPWR _0698_ _0772_ _0778_ _0779_ sky130_fd_sc_hd__o21a_1
X_6646_ VGND VPWR VPWR VGND _3035_ _3034_ _2993_ _3033_ sky130_fd_sc_hd__mux2_1
X_3858_ VGND VPWR VPWR VGND _0710_ _0670_ _0667_ i_tinyqv.cpu.i_core.i_registers.reg_access\[2\]\[0\]
+ net25 i_tinyqv.cpu.i_core.i_registers.reg_access\[8\]\[0\] sky130_fd_sc_hd__a32o_1
X_6577_ VPWR VGND VGND VPWR _2980_ _1400_ i_tinyqv.cpu.instr_data\[2\]\[0\] sky130_fd_sc_hd__or2_1
X_3789_ VPWR VGND VPWR VGND _0637_ i_tinyqv.cpu.i_core.i_registers.reg_access\[11\]\[3\]
+ _0640_ _0641_ sky130_fd_sc_hd__a21o_1
X_8316_ i_tinyqv.mem.q_ctrl.spi_in_buffer\[4\] clknet_leaf_18_clk _0415_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5528_ VPWR VGND VPWR VGND _2230_ net164 i_uart_tx.fsm_state\[3\] _2232_ sky130_fd_sc_hd__a21oi_1
X_5459_ VPWR VGND VGND VPWR _2184_ _2179_ _2183_ sky130_fd_sc_hd__or2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.i_regbuf\[12\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[12\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[16\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_8247_ i_tinyqv.cpu.i_core.mepc\[18\] clknet_leaf_34_clk _0347_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_8178_ i_tinyqv.cpu.instr_data\[1\]\[13\] clknet_leaf_13_clk _0290_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_580 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7129_ VPWR VGND VPWR VGND _3308_ _1483_ _2132_ _3435_ _2126_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_514 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_4830_ VGND VPWR _0038_ _1654_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4761_ VPWR VGND VGND VPWR _0894_ _1595_ _1596_ sky130_fd_sc_hd__nor2_1
X_6500_ VGND VPWR VGND VPWR _2914_ _2906_ i_tinyqv.mem.qspi_data_byte_idx\[1\] sky130_fd_sc_hd__xnor2_4
X_4692_ VGND VPWR _1527_ _1528_ _1526_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_7480_ VGND VPWR _3720_ i_tinyqv.cpu.instr_data_start\[20\] i_tinyqv.cpu.instr_data_start\[21\]
+ _3707_ VPWR VGND sky130_fd_sc_hd__and3_1
X_6431_ VPWR VGND VGND VPWR _2795_ _2864_ _2802_ sky130_fd_sc_hd__nand2_1
X_6362_ VPWR VGND _2795_ _2803_ _2802_ VPWR VGND sky130_fd_sc_hd__and2_2
X_8101_ i_tinyqv.cpu.instr_data\[1\]\[1\] clknet_leaf_9_clk _0213_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5313_ _2060_ _0707_ _0697_ _0814_ _2059_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
X_6293_ VGND VPWR VPWR VGND _2756_ _2322_ _1552_ net229 sky130_fd_sc_hd__mux2_1
X_5244_ VGND VPWR VPWR VGND _1995_ _0027_ _1997_ sky130_fd_sc_hd__xor2_1
X_8032_ i_tinyqv.cpu.instr_data\[3\]\[10\] clknet_leaf_4_clk _0167_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5175_ VGND VPWR _1904_ _1930_ _1931_ _1903_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_4126_ VPWR VGND _0973_ net28 _0907_ VPWR VGND sky130_fd_sc_hd__and2_1
X_4057_ VPWR VGND VPWR VGND _0888_ _0884_ i_tinyqv.cpu.instr_data_start\[4\] _0904_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_7816_ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[3\] clknet_leaf_1_clk _0073_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.i_regbuf\[24\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[24\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[28\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4959_ VGND VPWR _1735_ gpio_out\[4\] _1729_ _1730_ VPWR VGND sky130_fd_sc_hd__and3_1
X_7747_ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[30\] clknet_leaf_0_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[30\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_466 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7678_ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[25\] clknet_leaf_55_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[25\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6629_ VPWR VGND VPWR VGND i_tinyqv.cpu.i_core.imm_lo\[2\] net60 _2998_ _3022_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_171 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_14_160 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.i_regbuf\[13\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[13\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[17\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.i_regbuf\[8\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[8\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[12\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_200 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_52_288 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.i_regbuf\[12\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[12\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[16\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_cycles.i_regbuf\[10\] i_tinyqv.cpu.i_core.i_cycles.reg_buf\[10\]
+ i_tinyqv.cpu.i_core.i_cycles.register\[14\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6980_ VPWR VGND VPWR VGND _2119_ _3301_ _1483_ _3302_ sky130_fd_sc_hd__or3_1
X_5931_ VGND VPWR VPWR VGND _2519_ i_tinyqv.cpu.i_core.mepc\[8\] _2106_ i_tinyqv.cpu.i_core.i_shift.a\[12\]
+ sky130_fd_sc_hd__mux2_1
X_5862_ VGND VPWR _0219_ _2475_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5793_ VPWR VGND VPWR VGND _2339_ _2425_ _2198_ _2426_ sky130_fd_sc_hd__or3_1
X_4813_ VGND VPWR _0047_ _1644_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7601_ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[12\] clknet_leaf_0_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[12\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_583 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7532_ i_tinyqv.cpu.i_core.i_registers.reg_access\[15\]\[3\] clknet_leaf_45_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[7\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4744_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[2\] _1579_ _1250_ sky130_fd_sc_hd__nand2_1
X_7463_ VPWR VGND VPWR VGND i_tinyqv.mem.q_ctrl.addr\[14\] _2732_ _3706_ _3704_ _3705_
+ _3008_ sky130_fd_sc_hd__a221o_1
X_4675_ VPWR VGND VGND VPWR _1507_ _1511_ _1510_ sky130_fd_sc_hd__nand2_1
X_6414_ _2850_ _2803_ _2845_ _2847_ _2849_ _2837_ VPWR VGND VGND VPWR sky130_fd_sc_hd__o311a_1
X_7394_ VPWR VGND VPWR VGND _3648_ _2877_ _3647_ _3017_ _3080_ sky130_fd_sc_hd__a211oi_1
X_6345_ VPWR VGND VGND VPWR _2786_ _1707_ _2785_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_664 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_3_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_6276_ VGND VPWR _0361_ _2747_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8015_ i_uart_rx.bit_sample clknet_leaf_27_clk _0150_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5227_ VPWR VGND VGND VPWR _1978_ _1981_ _1980_ sky130_fd_sc_hd__nand2_1
X_5158_ VPWR VGND VGND VPWR _1913_ _1915_ _1914_ sky130_fd_sc_hd__nand2_1
X_4109_ VPWR VGND _0956_ _0688_ VPWR VGND sky130_fd_sc_hd__buf_2
X_5089_ VGND VPWR VGND VPWR _1848_ _1820_ _1821_ _1849_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_2_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_62_520 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_50_704 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_15_480 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.i_regbuf\[24\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[24\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[28\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_586 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_7_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_4460_ VGND VPWR VGND VPWR _1303_ _1243_ _1218_ _1302_ _1034_ _0877_ sky130_fd_sc_hd__a32o_2
X_4391_ VGND VPWR VGND VPWR _1234_ _1224_ _1230_ _0945_ _1233_ sky130_fd_sc_hd__o211a_1
X_6130_ VGND VPWR VPWR VGND _2639_ _2638_ _2468_ i_tinyqv.cpu.instr_data_in\[1\] sky130_fd_sc_hd__mux2_1
X_6061_ VGND VPWR _0295_ _2598_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5012_ VGND VPWR _1774_ _1775_ i_tinyqv.cpu.i_core.multiplier.accum\[4\] VPWR VGND
+ sky130_fd_sc_hd__xnor2_1
X_6963_ VGND VPWR VPWR VGND _3286_ i_tinyqv.cpu.instr_data\[2\]\[11\] _1504_ i_tinyqv.cpu.instr_data\[0\]\[11\]
+ sky130_fd_sc_hd__mux2_1
X_5914_ VGND VPWR VPWR VGND _2508_ _2507_ _2502_ i_tinyqv.cpu.data_addr\[2\] sky130_fd_sc_hd__mux2_1
X_6894_ VPWR VGND _3254_ _3253_ _0752_ VPWR VGND sky130_fd_sc_hd__and2_1
X_5845_ VPWR VGND VGND VPWR _2465_ _1400_ i_tinyqv.cpu.instr_data\[1\]\[1\] sky130_fd_sc_hd__or2_1
X_5776_ VGND VPWR VPWR VGND _2402_ _2404_ i_spi.bits_remaining\[2\] _2414_ sky130_fd_sc_hd__or3b_1
X_8564_ i_tinyqv.cpu.i_core.i_instrret.register\[3\] clknet_leaf_47_clk _0606_ VPWR
+ VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4727_ VGND VPWR VPWR VGND uo_out[7] _1549_ gpio_out_sel\[7\] _1561_ _1562_ sky130_fd_sc_hd__o31a_4
X_8495_ i_tinyqv.mem.q_ctrl.addr\[21\] clknet_leaf_32_clk _0593_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_2
X_7515_ VGND VPWR _0600_ _3747_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7446_ VPWR VGND VPWR VGND _3681_ _0881_ i_tinyqv.cpu.instr_data_start\[16\] _3691_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4658_ VPWR VGND VGND VPWR _1494_ _1452_ _1493_ sky130_fd_sc_hd__or2_1
X_7377_ VPWR VGND _3633_ i_tinyqv.cpu.instr_write_offset\[3\] _0884_ i_tinyqv.cpu.instr_data_start\[4\]
+ i_tinyqv.cpu.instr_data_start\[5\] VGND VPWR sky130_fd_sc_hd__a31o_1
X_4589_ VGND VPWR VGND VPWR _1425_ i_tinyqv.cpu.instr_data\[2\]\[1\] _1422_ _1408_
+ _1424_ sky130_fd_sc_hd__o211a_1
X_6328_ VGND VPWR _0385_ _2775_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6259_ VPWR VGND VGND VPWR i_tinyqv.mem.q_ctrl.data_ready i_tinyqv.mem.q_ctrl.data_req
+ _2735_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_634 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_39_325 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_11_Right_11 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Right_20 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_3960_ VPWR VGND VPWR VGND i_tinyqv.cpu.i_core.imm_lo\[2\] _0615_ _0812_ _0690_ i_tinyqv.cpu.i_core.imm_lo\[10\]
+ i_tinyqv.cpu.counter\[4\] sky130_fd_sc_hd__a221o_1
X_3891_ VPWR VGND VPWR VGND _0722_ _0721_ _0742_ _0743_ sky130_fd_sc_hd__a21o_1
X_5630_ VPWR VGND VGND VPWR _1543_ _2305_ _0158_ sky130_fd_sc_hd__nor2_1
X_5561_ VGND VPWR _2256_ i_uart_rx.cycle_counter\[8\] i_uart_rx.cycle_counter\[7\]
+ _2253_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_41_501 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5492_ VGND VPWR _2203_ _2200_ _2207_ net219 VPWR VGND sky130_fd_sc_hd__o21ai_1
X_8280_ i_tinyqv.mem.data_from_read\[20\] clknet_leaf_13_clk _0379_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_7300_ VPWR VGND VPWR VGND _3291_ _1486_ _3574_ _1510_ _3572_ _3573_ sky130_fd_sc_hd__a221o_1
X_4512_ VGND VPWR VPWR VGND _1351_ i_tinyqv.cpu.i_core.cycle_count_wide\[5\] _0841_
+ i_tinyqv.cpu.i_core.time_hi\[1\] sky130_fd_sc_hd__mux2_1
Xhold104 net133 i_tinyqv.mem.q_ctrl.spi_in_buffer\[1\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 VGND VPWR i_tinyqv.mem.q_ctrl.spi_clk_out net155 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xhold115 net144 i_tinyqv.cpu.load_started VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7231_ VPWR VGND _3519_ _3418_ _3330_ _3291_ _3510_ VGND VPWR sky130_fd_sc_hd__a31o_1
Xhold159 net188 i_debug_uart_tx.cycle_counter\[1\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 net166 _0130_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 net177 i_tinyqv.cpu.data_addr\[22\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_4443_ VGND VPWR VPWR VGND _1286_ _1130_ _1108_ _1127_ sky130_fd_sc_hd__mux2_1
X_7162_ VPWR VGND VGND VPWR _3368_ i_tinyqv.cpu.instr_data\[1\]\[15\] _3366_ i_tinyqv.cpu.instr_data\[0\]\[15\]
+ _3464_ _3463_ sky130_fd_sc_hd__o221a_2
X_4374_ VGND VPWR _0857_ _1216_ _1217_ _0777_ VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_6113_ VGND VPWR _2624_ _2625_ VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_7093_ VGND VPWR VPWR VGND _3403_ _3402_ _3319_ _2165_ sky130_fd_sc_hd__mux2_1
X_6044_ VGND VPWR VPWR VGND _2588_ i_tinyqv.cpu.instr_data\[1\]\[12\] _2462_ _1712_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7995_ i_uart_tx.fsm_state\[3\] clknet_leaf_30_clk net166 VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6946_ VGND VPWR VPWR VGND _0501_ _3274_ _3261_ _1589_ _3277_ net114 sky130_fd_sc_hd__a32o_1
XFILLER_0_49_623 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_6877_ VPWR VGND VGND VPWR i_tinyqv.cpu.is_store _3243_ _1761_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_14_Left_95 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_48_155 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5828_ VPWR VGND VPWR VGND _2088_ net66 _2434_ _2453_ sky130_fd_sc_hd__a21o_1
X_5759_ VGND VPWR VPWR VGND _2401_ i_spi.data\[0\] _2400_ _2391_ sky130_fd_sc_hd__mux2_1
X_8547_ i_tinyqv.cpu.i_core.i_cycles.register\[20\] clknet_leaf_51_clk i_tinyqv.cpu.i_core.i_cycles.reg_buf\[20\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_8478_ i_tinyqv.mem.q_ctrl.addr\[4\] clknet_leaf_29_clk _0576_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_7429_ VPWR VGND VGND VPWR i_tinyqv.cpu.was_early_branch _3676_ _3677_ sky130_fd_sc_hd__nor2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.i_regbuf\[27\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[27\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[31\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_38 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4090_ VGND VPWR VGND VPWR _0932_ i_tinyqv.cpu.i_core.imm_lo\[6\] _0937_ _0936_ sky130_fd_sc_hd__nand3_2
X_6800_ VPWR VGND VGND VPWR i_tinyqv.cpu.instr_data_start\[17\] _3175_ i_tinyqv.cpu.imm\[17\]
+ sky130_fd_sc_hd__nand2_1
X_7780_ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[31\] clknet_leaf_58_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[31\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4992_ VPWR VGND VPWR VGND _1754_ _1755_ _1604_ _1410_ _1756_ sky130_fd_sc_hd__or4_1
X_6731_ VGND VPWR VGND VPWR _0451_ i_tinyqv.cpu.instr_data_start\[10\] _3027_ _3112_
+ _3093_ sky130_fd_sc_hd__o211a_1
X_3943_ VPWR VGND VPWR VGND _0631_ i_tinyqv.cpu.i_core.i_registers.reg_access\[15\]\[2\]
+ _0633_ _0795_ i_tinyqv.cpu.i_core.i_registers.reg_access\[12\]\[2\] sky130_fd_sc_hd__a22o_1
X_6662_ VPWR VGND VGND VPWR _3037_ _3050_ _3049_ sky130_fd_sc_hd__nand2_1
X_3874_ VGND VPWR i_tinyqv.cpu.instr_data_start\[12\] _0726_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_5613_ VGND VPWR VGND VPWR _0153_ i_uart_rx.fsm_state\[1\] _2281_ _2293_ _2182_ sky130_fd_sc_hd__o211a_1
X_8401_ i_tinyqv.cpu.data_out\[26\] clknet_leaf_19_clk _0499_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_2__f_clk VGND VPWR VGND VPWR clknet_0_clk clknet_3_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_6593_ VPWR VGND _2991_ _2990_ VPWR VGND sky130_fd_sc_hd__buf_4
X_8332_ i_tinyqv.cpu.instr_data\[2\]\[1\] clknet_leaf_13_clk _0431_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5544_ VGND VPWR _2236_ _2242_ _2245_ net178 VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_60 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5475_ VGND VPWR VGND VPWR _0114_ net316 _2169_ _2194_ _2182_ sky130_fd_sc_hd__o211a_1
X_8263_ i_tinyqv.cpu.instr_data_in\[3\] clknet_leaf_14_clk _0362_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_14_589 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_30_93 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_8194_ i_tinyqv.cpu.i_core.i_shift.a\[13\] clknet_leaf_41_clk _0306_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
X_4426_ VPWR VGND VPWR VGND _1266_ _1092_ _1268_ _1269_ sky130_fd_sc_hd__a21oi_1
X_7214_ VPWR VGND _3508_ _3507_ _3476_ _3328_ _3362_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_7145_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.imm_lo\[8\] _3360_ _3449_ _0528_ sky130_fd_sc_hd__o21a_1
X_4357_ VPWR VGND VPWR VGND _0894_ _0726_ i_tinyqv.cpu.instr_data_start\[13\] _1200_
+ sky130_fd_sc_hd__a21oi_1
X_4288_ VGND VPWR VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[25\] i_tinyqv.cpu.i_core.i_shift.a\[26\]
+ i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt\[0\] i_tinyqv.cpu.i_core.i_shift.a\[6\]
+ i_tinyqv.cpu.i_core.i_shift.a\[5\] _1029_ _1135_ sky130_fd_sc_hd__mux4_1
X_7076_ VGND VPWR _0521_ _3387_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6027_ VGND VPWR _0280_ _2579_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7978_ i_uart_tx.data_to_send\[5\] clknet_leaf_28_clk _0113_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_6929_ VPWR VGND VPWR VGND _3272_ _3253_ _3261_ _0489_ net156 sky130_fd_sc_hd__a22o_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.i_regbuf\[28\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[28\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5260_ VPWR VGND VGND VPWR _2011_ _2013_ _2012_ sky130_fd_sc_hd__nand2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.i_regbuf\[31\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[31\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[3\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4211_ VPWR VGND _1042_ _1058_ _1057_ VPWR VGND sky130_fd_sc_hd__and2_2
X_5191_ VPWR VGND _1947_ _1946_ _1945_ VPWR VGND sky130_fd_sc_hd__and2_1
X_4142_ VGND VPWR VGND VPWR _0988_ i_debug_uart_tx.fsm_state\[0\] _0989_ sky130_fd_sc_hd__or2_4
X_4073_ VPWR VGND VGND VPWR _0919_ _0920_ _0855_ sky130_fd_sc_hd__nor2_2
X_7901_ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[24\] clknet_leaf_48_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[24\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_559 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_7832_ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[19\] clknet_leaf_52_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[19\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4975_ VGND VPWR _1745_ gpio_out_sel\[2\] _1737_ _1742_ VPWR VGND sky130_fd_sc_hd__and3_1
X_7763_ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[14\] clknet_leaf_53_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[14\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_401 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6714_ VPWR VGND VGND VPWR _3097_ _0882_ i_tinyqv.cpu.i_core.imm_lo\[9\] sky130_fd_sc_hd__or2_1
XFILLER_0_19_648 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_3926_ VPWR VGND VGND VPWR _0698_ _0778_ _0777_ sky130_fd_sc_hd__nand2_1
X_7694_ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[9\] clknet_leaf_53_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[9\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_659 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_6645_ VGND VPWR VPWR VGND _3034_ _3023_ _2991_ _2509_ sky130_fd_sc_hd__mux2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.i_regbuf\[16\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[16\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[20\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3857_ VPWR VGND VPWR VGND net24 i_tinyqv.cpu.i_core.i_registers.reg_access\[15\]\[0\]
+ _0677_ _0709_ i_tinyqv.cpu.i_core.i_registers.reg_access\[1\]\[0\] sky130_fd_sc_hd__a22o_1
X_6576_ VPWR VGND VGND VPWR _2229_ _1543_ _0429_ sky130_fd_sc_hd__nor2_1
X_3788_ VPWR VGND VPWR VGND _0639_ i_tinyqv.cpu.i_core.i_registers.reg_access\[2\]\[3\]
+ _0638_ _0640_ i_tinyqv.cpu.i_core.i_registers.reg_access\[6\]\[3\] sky130_fd_sc_hd__a22o_1
X_8315_ i_tinyqv.mem.q_ctrl.spi_in_buffer\[3\] clknet_leaf_16_clk _0414_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5527_ VPWR VGND VGND VPWR _2229_ _2231_ _0129_ sky130_fd_sc_hd__nor2_1
X_8246_ i_tinyqv.cpu.i_core.mepc\[17\] clknet_leaf_35_clk _0346_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_5458_ VGND VPWR VPWR VGND _2183_ i_uart_tx.data_to_send\[2\] _2177_ i_uart_tx.data_to_send\[1\]
+ sky130_fd_sc_hd__mux2_1
X_4409_ VGND VPWR VPWR VGND _1249_ _1252_ _1251_ sky130_fd_sc_hd__xor2_1
X_5389_ VPWR VGND VGND VPWR _2119_ _1469_ _2118_ sky130_fd_sc_hd__or2_1
X_8177_ i_tinyqv.cpu.instr_data\[1\]\[12\] clknet_leaf_10_clk _0289_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_7128_ VPWR VGND VGND VPWR _3368_ i_tinyqv.cpu.instr_data\[1\]\[11\] _3366_ i_tinyqv.cpu.instr_data\[0\]\[11\]
+ _3434_ _3433_ sky130_fd_sc_hd__o221a_1
X_7059_ VGND VPWR _3371_ _3372_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_65_710 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_37_445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_33_640 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_20_345 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_412 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4760_ VPWR VGND VGND VPWR i_tinyqv.cpu.instr_data_start\[11\] _0893_ _1595_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_445 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4691_ VGND VPWR _1522_ _1527_ i_tinyqv.cpu.instr_write_offset\[3\] VPWR VGND sky130_fd_sc_hd__xnor2_1
X_6430_ VGND VPWR VGND VPWR _2863_ _2860_ _2836_ _2862_ _2806_ sky130_fd_sc_hd__o211a_1
X_6361_ VPWR VGND VGND VPWR i_tinyqv.mem.q_ctrl.delay_cycles_cfg\[2\] _2802_ _2789_
+ sky130_fd_sc_hd__nand2_1
X_8100_ i_tinyqv.cpu.instr_data\[1\]\[0\] clknet_leaf_8_clk _0212_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_49_Right_49 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5312_ VPWR VGND VGND VPWR _0777_ _2055_ _2059_ sky130_fd_sc_hd__nor2_1
X_6292_ VGND VPWR _0369_ _2755_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5243_ VPWR VGND VGND VPWR _1969_ _1997_ _1996_ sky130_fd_sc_hd__nand2_1
X_8031_ i_tinyqv.cpu.instr_data\[3\]\[9\] clknet_leaf_10_clk _0166_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5174_ VPWR VGND VGND VPWR _1930_ _1929_ _1924_ sky130_fd_sc_hd__or2_1
X_4125_ VPWR VGND VGND VPWR i_tinyqv.cpu.data_addr\[25\] i_tinyqv.cpu.data_addr\[26\]
+ i_tinyqv.cpu.data_addr\[27\] _0972_ sky130_fd_sc_hd__nor3_1
XPHY_EDGE_ROW_58_Right_58 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4056_ VPWR VGND VGND VPWR _0610_ _0903_ _0902_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7815_ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[2\] clknet_leaf_57_clk _0072_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4958_ VPWR VGND VPWR VGND _1727_ net197 _1734_ _0003_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_551 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7746_ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[29\] clknet_leaf_55_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[29\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_434 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.i_regbuf\[17\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[17\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[21\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7677_ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[24\] clknet_leaf_59_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[24\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_3909_ VGND VPWR VGND VPWR _0761_ net63 _0758_ i_tinyqv.cpu.i_core.i_registers.reg_access\[13\]\[1\]
+ _0760_ sky130_fd_sc_hd__a211o_1
X_4889_ VGND VPWR VPWR VGND _1688_ _1380_ _1685_ i_tinyqv.cpu.i_core.i_registers.reg_access\[6\]\[2\]
+ sky130_fd_sc_hd__mux2_1
X_6628_ VPWR VGND VGND VPWR _3019_ _3021_ _3020_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_67_Right_67 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6559_ VPWR VGND VGND VPWR _2967_ i_tinyqv.cpu.data_out\[30\] _2912_ sky130_fd_sc_hd__or2_1
X_8229_ i_tinyqv.cpu.i_core.mepc\[0\] clknet_leaf_35_clk _0329_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_76_Right_76 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.i_regbuf\[20\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[20\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[24\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_710 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_25_459 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_2_Left_83 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.i_regbuf\[8\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[8\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[12\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_643 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_5930_ VGND VPWR _0244_ _2518_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7600_ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[11\] clknet_leaf_1_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[11\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5861_ VGND VPWR VPWR VGND _2475_ i_tinyqv.cpu.instr_data\[0\]\[7\] _2469_ i_tinyqv.cpu.instr_data_in\[7\]
+ sky130_fd_sc_hd__mux2_1
X_5792_ VPWR VGND VGND VPWR net205 _2334_ _0988_ _2425_ sky130_fd_sc_hd__o21a_1
X_4812_ VGND VPWR VPWR VGND _1644_ i_tinyqv.cpu.debug_rd\[1\] _1642_ i_tinyqv.cpu.i_core.i_registers.reg_access\[14\]\[1\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_659 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_7531_ i_tinyqv.cpu.i_core.i_registers.reg_access\[15\]\[2\] clknet_leaf_44_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[6\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4743_ VGND VPWR _1578_ _1570_ _1577_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_7462_ VPWR VGND VGND VPWR i_tinyqv.cpu.data_addr\[18\] _2681_ _3004_ _3705_ sky130_fd_sc_hd__o21a_1
XFILLER_0_7_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_22_72 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6413_ VPWR VGND VPWR VGND i_tinyqv.mem.q_ctrl.nibbles_remaining\[0\] i_tinyqv.mem.q_ctrl.nibbles_remaining\[1\]
+ _2848_ _2849_ sky130_fd_sc_hd__a21o_1
X_4674_ VGND VPWR VPWR VGND _1510_ _1432_ _1509_ _1508_ sky130_fd_sc_hd__mux2_4
X_7393_ VPWR VGND VGND VPWR _3645_ _3646_ _3239_ _3647_ sky130_fd_sc_hd__o21a_1
X_6344_ VPWR VGND VGND VPWR _1706_ _2785_ i_tinyqv.mem.q_ctrl.fsm_state\[1\] sky130_fd_sc_hd__nand2_1
X_6275_ VGND VPWR VPWR VGND _2747_ i_tinyqv.cpu.instr_data_in\[2\] _2744_ _2320_ sky130_fd_sc_hd__mux2_1
X_8014_ i_uart_rx.recieved_data\[7\] clknet_leaf_28_clk _0149_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5226_ VGND VPWR _1953_ _1979_ _1980_ _1952_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_5157_ VPWR VGND VGND VPWR _1901_ _1887_ _1914_ _1912_ sky130_fd_sc_hd__nand3_1
X_4108_ VGND VPWR VGND VPWR _0955_ _0752_ i_tinyqv.cpu.i_core.mem_op\[0\] _0945_ i_tinyqv.cpu.i_core.mem_op\[1\]
+ sky130_fd_sc_hd__a211o_2
X_5088_ _1848_ _1817_ _1819_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.i_regbuf\[7\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[7\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[11\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4039_ VPWR VGND VGND VPWR i_tinyqv.cpu.instr_len\[2\] i_tinyqv.cpu.pc\[2\] _0886_
+ sky130_fd_sc_hd__nor2_1
X_7729_ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[12\] clknet_leaf_59_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[12\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_584 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_6_191 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.i_regbuf\[21\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[21\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[25\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.i_regbuf\[10\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[10\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[14\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.i_regbuf\[17\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[17\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[21\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_40_215 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_4390_ VGND VPWR VGND VPWR _1233_ net14 _1231_ gpio_out_sel\[5\] _1232_ sky130_fd_sc_hd__a211o_1
X_6060_ VGND VPWR VPWR VGND _2598_ i_tinyqv.cpu.i_core.i_shift.a\[2\] _2596_ i_tinyqv.cpu.i_core.i_shift.a\[6\]
+ sky130_fd_sc_hd__mux2_1
X_5011_ VGND VPWR VPWR VGND _1771_ _1774_ _1773_ sky130_fd_sc_hd__xor2_1
X_6962_ VGND VPWR VPWR VGND _3285_ i_tinyqv.cpu.instr_data\[3\]\[11\] _1504_ i_tinyqv.cpu.instr_data\[1\]\[11\]
+ sky130_fd_sc_hd__mux2_1
X_6893_ VPWR VGND VGND VPWR _0854_ _3253_ _0612_ sky130_fd_sc_hd__nor2_2
X_5913_ VGND VPWR VPWR VGND _2504_ i_tinyqv.cpu.i_core.mepc\[2\] i_tinyqv.cpu.i_core.i_shift.a\[6\]
+ _2507_ sky130_fd_sc_hd__mux2_2
X_5844_ VGND VPWR _0212_ _2464_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8563_ i_tinyqv.cpu.i_core.i_instrret.register\[2\] clknet_leaf_50_clk _0605_ VPWR
+ VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5775_ VGND VPWR _0195_ _2413_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7514_ VGND VPWR _3747_ net90 _1752_ _3746_ VPWR VGND sky130_fd_sc_hd__and3_1
X_4726_ VGND VPWR VGND VPWR gpio_out\[7\] _1562_ gpio_out_sel\[7\] sky130_fd_sc_hd__or2b_1
X_8494_ i_tinyqv.mem.q_ctrl.addr\[20\] clknet_leaf_32_clk _0592_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_2
X_7445_ VGND VPWR _3690_ _0881_ i_tinyqv.cpu.instr_data_start\[16\] _3681_ VPWR VGND
+ sky130_fd_sc_hd__and3_1
X_4657_ VPWR VGND VPWR VGND _1491_ _1492_ _1455_ _1493_ sky130_fd_sc_hd__or3_4
X_7376_ VGND VPWR i_tinyqv.cpu.was_early_branch _3632_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_6327_ VGND VPWR VPWR VGND _2775_ _2320_ _2772_ net267 sky130_fd_sc_hd__mux2_1
X_4588_ VPWR VGND VGND VPWR _1424_ i_tinyqv.cpu.instr_data\[0\]\[1\] net36 sky130_fd_sc_hd__or2_1
X_6258_ VPWR VGND VGND VPWR _2679_ _2734_ i_tinyqv.mem.instr_active sky130_fd_sc_hd__nor2_2
X_5209_ VPWR VGND VGND VPWR _1932_ _1935_ _1964_ _1962_ sky130_fd_sc_hd__nand3_1
X_6189_ VGND VPWR _0346_ _2675_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_576 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_3890_ VGND VPWR VPWR VGND _0742_ _0654_ _0741_ _0729_ sky130_fd_sc_hd__mux2_4
X_5560_ VPWR VGND VPWR VGND _2253_ net199 _2255_ _0138_ sky130_fd_sc_hd__a21oi_1
X_5491_ VPWR VGND _2206_ _2203_ i_uart_tx.cycle_counter\[3\] VPWR VGND sky130_fd_sc_hd__and2_1
X_4511_ VPWR VGND VPWR VGND _0841_ _0946_ _0934_ _1350_ sky130_fd_sc_hd__a21oi_1
Xhold105 net134 _2903_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 net145 i_tinyqv.mem.q_ctrl.spi_data_oe\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7230_ VGND VPWR _0544_ _3518_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4442_ VGND VPWR VPWR VGND _1285_ _1126_ _1108_ _1155_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_557 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold149 net178 i_uart_rx.cycle_counter\[2\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 net167 i_tinyqv.mem.q_ctrl.spi_in_buffer\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 net156 i_tinyqv.cpu.data_out\[16\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7161_ VPWR VGND VPWR VGND i_tinyqv.cpu.instr_data\[3\]\[15\] _3369_ _3463_ _3370_
+ i_tinyqv.cpu.instr_data\[2\]\[15\] _3372_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_4373_ VGND VPWR VGND VPWR _1216_ _1199_ _1215_ _0921_ _0880_ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6112_ VPWR VGND VGND VPWR _2624_ _0846_ _1755_ sky130_fd_sc_hd__or2_1
X_7092_ VPWR VGND VGND VPWR _3368_ i_tinyqv.cpu.instr_data\[1\]\[7\] _3366_ i_tinyqv.cpu.instr_data\[0\]\[7\]
+ _3402_ _3401_ sky130_fd_sc_hd__o221a_1
X_6043_ VGND VPWR _0288_ _2587_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_71 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_7994_ i_uart_tx.fsm_state\[2\] clknet_leaf_29_clk _0129_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_14_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6945_ VPWR VGND VGND VPWR _3277_ _1604_ _0854_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_635 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_6876_ VPWR VGND _0466_ _1604_ _2049_ _3017_ _1480_ VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_76_498 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_5827_ VPWR VGND VPWR VGND _2452_ _2451_ _2083_ _0208_ sky130_fd_sc_hd__a21oi_1
X_5758_ VPWR VGND VPWR VGND _2397_ i_spi.read_latency _2399_ _2400_ sky130_fd_sc_hd__a21oi_1
X_8546_ i_tinyqv.cpu.i_core.i_cycles.register\[19\] clknet_leaf_50_clk i_tinyqv.cpu.i_core.i_cycles.reg_buf\[19\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4709_ VGND VPWR VGND VPWR net5 _1543_ _1532_ _1544_ _0946_ _1385_ _1545_ sky130_fd_sc_hd__mux4_2
X_8477_ i_tinyqv.cpu.instr_write_offset\[3\] clknet_leaf_22_clk _0575_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_17_576 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5689_ VPWR VGND _2347_ _2337_ i_debug_uart_tx.data_to_send\[4\] VPWR VGND sky130_fd_sc_hd__and2_1
X_7428_ VGND VPWR _3676_ _0726_ i_tinyqv.cpu.instr_data_start\[13\] _3667_ VPWR VGND
+ sky130_fd_sc_hd__and3_1
X_7359_ VGND VPWR _1443_ _2147_ _3619_ _2993_ VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_307 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_6730_ VPWR VGND VGND VPWR _3037_ _3112_ _3111_ sky130_fd_sc_hd__nand2_1
X_4991_ VPWR VGND VPWR VGND _1755_ i_tinyqv.cpu.i_core.cycle\[1\] i_tinyqv.cpu.i_core.cycle\[0\]
+ sky130_fd_sc_hd__or2_2
X_3942_ VPWR VGND VPWR VGND net26 i_tinyqv.cpu.i_core.i_registers.reg_access\[8\]\[2\]
+ net27 _0794_ i_tinyqv.cpu.i_core.i_registers.reg_access\[2\]\[2\] sky130_fd_sc_hd__a22o_1
X_6661_ VPWR VGND VPWR VGND _3038_ _3039_ _3049_ _2995_ _0905_ _3048_ sky130_fd_sc_hd__a221o_1
X_3873_ VPWR VGND VGND VPWR i_tinyqv.cpu.counter\[4\] _0724_ _0725_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_318 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5612_ VGND VPWR VGND VPWR _2292_ _2291_ _2289_ _1227_ _2290_ _2293_ sky130_fd_sc_hd__a311o_1
X_8400_ i_tinyqv.cpu.data_out\[25\] clknet_leaf_26_clk _0498_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_6592_ VGND VPWR _2989_ _2990_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_5543_ VPWR VGND VGND VPWR _2236_ _2244_ _0132_ sky130_fd_sc_hd__nor2_1
X_8331_ i_tinyqv.cpu.instr_data\[2\]\[0\] clknet_leaf_13_clk _0430_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5474_ VPWR VGND VGND VPWR _2194_ _2179_ _2193_ sky130_fd_sc_hd__or2_1
X_8262_ i_tinyqv.cpu.instr_data_in\[2\] clknet_leaf_14_clk _0361_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_7213_ VPWR VGND VPWR VGND i_tinyqv.cpu.instr_data\[0\]\[3\] _3487_ _3507_ _3488_
+ i_tinyqv.cpu.instr_data\[1\]\[3\] _3506_ sky130_fd_sc_hd__a221o_1
X_8193_ i_tinyqv.cpu.i_core.i_shift.a\[12\] clknet_leaf_41_clk _0305_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
X_4425_ VPWR VGND VPWR VGND _1267_ _1080_ _1077_ _1268_ sky130_fd_sc_hd__a21o_1
X_4356_ VGND VPWR VGND VPWR _1199_ net19 _1195_ i_tinyqv.cpu.i_core.mepc\[1\] _1198_
+ sky130_fd_sc_hd__a211o_1
X_7144_ VPWR VGND VPWR VGND _3443_ _3448_ _3362_ _3449_ sky130_fd_sc_hd__or3_1
X_4287_ VGND VPWR VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[3\] i_tinyqv.cpu.i_core.i_shift.a\[28\]
+ _1029_ i_tinyqv.cpu.i_core.i_shift.a\[4\] i_tinyqv.cpu.i_core.i_shift.a\[27\] _1103_
+ _1134_ sky130_fd_sc_hd__mux4_1
X_7075_ VGND VPWR VPWR VGND _3387_ _3386_ _3359_ i_tinyqv.cpu.i_core.imm_lo\[1\] sky130_fd_sc_hd__mux2_1
X_6026_ VGND VPWR VPWR VGND _2579_ i_tinyqv.cpu.instr_data\[1\]\[3\] _2463_ i_tinyqv.cpu.instr_data_in\[3\]
+ sky130_fd_sc_hd__mux2_1
X_7977_ i_uart_tx.data_to_send\[4\] clknet_leaf_28_clk _0112_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_6928_ VPWR VGND VGND VPWR _3272_ _0916_ _0854_ sky130_fd_sc_hd__or2_1
X_6859_ VGND VPWR VPWR VGND _3229_ _3228_ _2990_ _2548_ sky130_fd_sc_hd__mux2_1
X_8529_ i_tinyqv.cpu.i_core.i_cycles.register\[3\] clknet_leaf_51_clk _0599_ VPWR
+ VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_693 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_3_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_107 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_35_192 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_11_505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_387 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4210_ VPWR VGND VGND VPWR _1057_ i_tinyqv.cpu.i_core.i_shift.b\[2\] _1041_ sky130_fd_sc_hd__or2_1
X_5190_ VPWR VGND VGND VPWR _1946_ _1942_ _1943_ sky130_fd_sc_hd__or2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.i_regbuf\[24\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[24\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[28\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4141_ VGND VPWR VPWR VGND i_debug_uart_tx.fsm_state\[2\] i_debug_uart_tx.fsm_state\[1\]
+ i_debug_uart_tx.fsm_state\[3\] _0988_ sky130_fd_sc_hd__or3_2
X_4072_ VPWR VGND VGND VPWR i_tinyqv.cpu.alu_op\[0\] _0919_ _0656_ sky130_fd_sc_hd__nor2_2
X_7900_ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[23\] clknet_leaf_47_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[23\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7831_ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[18\] clknet_leaf_3_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[18\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4974_ VPWR VGND VPWR VGND _1741_ net97 _1744_ _0009_ sky130_fd_sc_hd__a21o_1
X_7762_ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[13\] clknet_leaf_54_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[13\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6713_ VPWR VGND VGND VPWR _0882_ _3096_ i_tinyqv.cpu.i_core.imm_lo\[9\] sky130_fd_sc_hd__nand2_1
X_3925_ VGND VPWR VGND VPWR _0611_ _0773_ _0776_ _0774_ _0777_ sky130_fd_sc_hd__o22a_2
X_7693_ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[8\] clknet_leaf_2_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[8\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6644_ VGND VPWR VPWR VGND _3033_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[11\]
+ net31 _1591_ sky130_fd_sc_hd__mux2_1
X_3856_ VPWR VGND VGND VPWR _0707_ _0708_ _0702_ sky130_fd_sc_hd__nor2_2
X_6575_ VGND VPWR _0428_ _2979_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_3787_ VGND VPWR VGND VPWR _0627_ _0639_ _0625_ _0624_ _0626_ sky130_fd_sc_hd__and4bb_2
X_8314_ i_tinyqv.mem.q_ctrl.spi_in_buffer\[2\] clknet_leaf_16_clk _0413_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5526_ VGND VPWR _2230_ _2231_ i_uart_tx.fsm_state\[2\] VPWR VGND sky130_fd_sc_hd__xnor2_1
X_5457_ VGND VPWR VGND VPWR _0108_ net117 _2169_ _2180_ _2182_ sky130_fd_sc_hd__o211a_1
X_8245_ i_tinyqv.cpu.i_core.mepc\[16\] clknet_leaf_35_clk _0345_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_4408_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[0\] _1251_ _1250_ sky130_fd_sc_hd__nand2_1
X_8176_ i_tinyqv.cpu.instr_data\[1\]\[11\] clknet_leaf_11_clk _0288_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5388_ VPWR VGND VPWR VGND _2118_ _1486_ sky130_fd_sc_hd__inv_2
X_7127_ VPWR VGND VPWR VGND i_tinyqv.cpu.instr_data\[3\]\[11\] _3369_ _3433_ _3370_
+ i_tinyqv.cpu.instr_data\[2\]\[11\] _3372_ sky130_fd_sc_hd__a221o_1
X_4339_ VPWR VGND VGND VPWR _1185_ _0855_ _0919_ sky130_fd_sc_hd__or2_1
X_7058_ VPWR VGND VGND VPWR _3365_ _3371_ _3367_ sky130_fd_sc_hd__nand2_1
X_6009_ VGND VPWR _0271_ _2570_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xi_tinyqv.cpu.i_core.i_cycles.i_regbuf\[7\] i_tinyqv.cpu.i_core.i_cycles.reg_buf\[7\]
+ i_tinyqv.cpu.i_core.i_cycles.register\[11\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_696 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_57_clk VGND VPWR clknet_3_0__leaf_clk clknet_leaf_57_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_4690_ VGND VPWR VPWR VGND _1440_ _0888_ _1439_ _1526_ sky130_fd_sc_hd__or3b_1
X_6360_ VPWR VGND VPWR VGND _2801_ _2800_ _2783_ sky130_fd_sc_hd__or2_2
XFILLER_0_70_257 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_51_471 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5311_ VGND VPWR VGND VPWR _2057_ _0922_ _2055_ _2058_ i_tinyqv.cpu.i_core.mcause\[0\]
+ sky130_fd_sc_hd__a2bb2o_1
X_6291_ VGND VPWR VPWR VGND _2755_ _2320_ _1552_ i_tinyqv.mem.qspi_data_buf\[10\]
+ sky130_fd_sc_hd__mux2_1
X_8030_ i_tinyqv.cpu.instr_data\[3\]\[8\] clknet_leaf_11_clk _0165_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.i_regbuf\[25\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[25\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[29\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5242_ VGND VPWR VGND VPWR _1996_ _1972_ _1945_ _1971_ sky130_fd_sc_hd__a21bo_1
X_5173_ VPWR VGND VGND VPWR _1054_ _1929_ _1880_ sky130_fd_sc_hd__nand2_1
X_4124_ VGND VPWR VGND VPWR _0969_ _0968_ _0970_ _0971_ sky130_fd_sc_hd__a21o_2
Xinput1 VPWR VGND net1 rst_n VPWR VGND sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_48_clk VGND VPWR clknet_3_4__leaf_clk clknet_leaf_48_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_4055_ VPWR VGND VGND VPWR _0900_ _0901_ _0902_ sky130_fd_sc_hd__nor2_1
X_7814_ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[1\] clknet_leaf_56_clk _0071_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4957_ VGND VPWR _1734_ gpio_out\[3\] _1729_ _1730_ VPWR VGND sky130_fd_sc_hd__and3_1
X_7745_ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[28\] clknet_leaf_0_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[28\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_457 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7676_ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[23\] clknet_leaf_46_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[23\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_3908_ VPWR VGND VPWR VGND i_tinyqv.cpu.i_core.i_registers.reg_access\[15\]\[1\]
+ net83 _0760_ net54 i_tinyqv.cpu.i_core.i_registers.reg_access\[9\]\[1\] _0759_ sky130_fd_sc_hd__a221o_1
X_4888_ VGND VPWR _0067_ _1687_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6627_ VPWR VGND VGND VPWR _3020_ i_tinyqv.cpu.instr_data_start\[3\] i_tinyqv.cpu.i_core.imm_lo\[3\]
+ sky130_fd_sc_hd__or2_1
X_3839_ VGND VPWR _0690_ _0691_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_34_438 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_6558_ VGND VPWR VPWR VGND _2966_ i_tinyqv.cpu.data_out\[14\] _2909_ i_debug_uart_tx.uart_tx_data\[6\]
+ sky130_fd_sc_hd__mux2_1
X_6489_ VGND VPWR _0417_ _2904_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5509_ VPWR VGND _2218_ _2215_ i_uart_tx.cycle_counter\[9\] VPWR VGND sky130_fd_sc_hd__and2_1
X_8228_ i_tinyqv.cpu.i_core.multiplier.accum\[11\] clknet_leaf_43_clk _0018_ VPWR
+ VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_8159_ i_tinyqv.cpu.instr_data\[2\]\[8\] clknet_leaf_11_clk _0271_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.i_regbuf\[13\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[13\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[17\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_39_clk VGND VPWR clknet_3_5__leaf_clk clknet_leaf_39_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_0_37_287 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_471 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_instrret.i_regbuf\[12\] i_tinyqv.cpu.i_core.i_instrret.reg_buf\[12\]
+ i_tinyqv.cpu.i_core.i_instrret.register\[16\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5860_ VGND VPWR _0218_ _2474_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4811_ VGND VPWR _0046_ _1643_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5791_ VGND VPWR _0200_ _2424_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7530_ i_tinyqv.cpu.i_core.i_registers.reg_access\[15\]\[1\] clknet_leaf_46_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[5\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4742_ VPWR VGND _1577_ _1576_ i_tinyqv.cpu.i_core.multiplier.accum\[3\] VPWR VGND
+ sky130_fd_sc_hd__xor2_2
X_7461_ VPWR VGND VGND VPWR _3012_ _3704_ _3703_ sky130_fd_sc_hd__nand2_1
X_4673_ VGND VPWR VPWR VGND _1509_ i_tinyqv.cpu.instr_data\[2\]\[7\] _1449_ i_tinyqv.cpu.instr_data\[0\]\[7\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_235 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_6412_ VGND VPWR i_tinyqv.mem.q_ctrl.nibbles_remaining\[0\] _2802_ _2848_ i_tinyqv.mem.q_ctrl.nibbles_remaining\[1\]
+ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_7392_ VPWR VGND VPWR VGND _3634_ _0883_ i_tinyqv.cpu.instr_data_start\[7\] _3646_
+ sky130_fd_sc_hd__a21oi_1
X_6343_ VPWR VGND VGND VPWR _2782_ _2783_ _2784_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_365 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6274_ VGND VPWR _0360_ _2746_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8013_ i_uart_rx.recieved_data\[6\] clknet_leaf_19_clk _0148_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_5225_ VPWR VGND VGND VPWR _1979_ _1925_ _1974_ sky130_fd_sc_hd__or2_1
X_5156_ VPWR VGND VPWR VGND _1887_ _1901_ _1912_ _1913_ sky130_fd_sc_hd__a21o_1
X_5087_ VGND VPWR VPWR VGND _1844_ _1847_ _1846_ sky130_fd_sc_hd__xor2_1
X_4107_ VPWR VGND VGND VPWR _0878_ _0954_ _0953_ sky130_fd_sc_hd__nand2_1
X_4038_ VPWR VGND _0885_ i_tinyqv.cpu.pc\[2\] i_tinyqv.cpu.instr_len\[2\] VPWR VGND
+ sky130_fd_sc_hd__and2_1
XFILLER_0_78_176 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_66_338 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5989_ VGND VPWR _0263_ _2558_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7728_ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[11\] clknet_leaf_53_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[11\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_298 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_7659_ i_tinyqv.cpu.i_core.i_registers.reg_access\[11\]\[2\] clknet_leaf_58_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[6\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.i_regbuf\[25\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[25\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[29\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.i_regbuf\[14\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[14\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[18\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_500 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_25_257 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5010_ VGND VPWR _1574_ _1772_ _1773_ _1573_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_6961_ VPWR VGND VPWR VGND _3284_ _3283_ sky130_fd_sc_hd__inv_2
X_5912_ VGND VPWR _0238_ _2506_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6892_ VPWR VGND _0472_ _1442_ net144 i_tinyqv.cpu.is_load _1760_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_5843_ VGND VPWR VPWR VGND _2464_ _2459_ _2463_ i_tinyqv.cpu.instr_data_in\[0\] sky130_fd_sc_hd__mux2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.i_regbuf\[5\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[5\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[9\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_8562_ i_tinyqv.cpu.i_core.i_instrret.register\[1\] clknet_leaf_48_clk _0604_ VPWR
+ VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5774_ VPWR VGND _2413_ _2412_ _2181_ VPWR VGND sky130_fd_sc_hd__and2_1
X_7513_ VPWR VGND _3746_ _3745_ i_tinyqv.cpu.i_core.i_instrret.data\[2\] VPWR VGND
+ sky130_fd_sc_hd__and2_1
XFILLER_0_29_596 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_4725_ VPWR VGND VPWR VGND _1554_ net7 _1560_ _1561_ sky130_fd_sc_hd__a21oi_1
X_8493_ i_tinyqv.mem.q_ctrl.addr\[19\] clknet_leaf_32_clk _0591_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_7444_ VPWR VGND VPWR VGND net303 _3007_ _0587_ _3009_ net318 _3689_ sky130_fd_sc_hd__a221o_1
X_4656_ VPWR VGND VGND VPWR _1492_ _1448_ _1460_ sky130_fd_sc_hd__or2_1
X_7375_ VPWR VGND VGND VPWR _3631_ _3625_ net151 _3630_ _0576_ sky130_fd_sc_hd__o22a_1
X_4587_ VPWR VGND VPWR VGND _1423_ i_tinyqv.cpu.instr_data\[3\]\[1\] _1422_ sky130_fd_sc_hd__or2_2
XFILLER_0_4_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_6326_ VGND VPWR _0384_ _2774_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6257_ VGND VPWR _2732_ _2733_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_5208_ VPWR VGND VPWR VGND _1935_ _1932_ _1962_ _1963_ sky130_fd_sc_hd__a21o_1
X_6188_ VGND VPWR VPWR VGND _2675_ i_tinyqv.cpu.i_core.mepc\[21\] _2667_ i_tinyqv.cpu.i_core.mepc\[17\]
+ sky130_fd_sc_hd__mux2_1
X_5139_ VPWR VGND VGND VPWR _1894_ _1897_ _1896_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_26_Left_107 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Left_116 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_26_522 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_5490_ VGND VPWR _0118_ _2205_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4510_ VPWR VGND VGND VPWR _0946_ _1348_ _1349_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold106 net135 i_tinyqv.cpu.imm\[31\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4441_ VGND VPWR VPWR VGND _1284_ _1283_ _1058_ _1282_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_44_Left_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold117 net146 i_tinyqv.cpu.imm\[29\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 net168 _2902_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold128 net157 i_uart_tx.cycle_counter\[7\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7160_ VGND VPWR _0530_ _3462_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_9_Right_9 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6111_ VGND VPWR _0320_ _2623_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4372_ VPWR VGND VPWR VGND _1214_ _1210_ _0858_ _1215_ sky130_fd_sc_hd__a21oi_1
X_7091_ VPWR VGND VPWR VGND i_tinyqv.cpu.instr_data\[3\]\[7\] _3369_ _3401_ _3370_
+ i_tinyqv.cpu.instr_data\[2\]\[7\] _3372_ sky130_fd_sc_hd__a221o_1
X_6042_ VGND VPWR VPWR VGND _2587_ i_tinyqv.cpu.instr_data\[1\]\[11\] _2462_ _2322_
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_53_Left_134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7993_ i_uart_tx.fsm_state\[1\] clknet_leaf_29_clk _0128_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6944_ VGND VPWR VPWR VGND _0500_ _3274_ _3269_ _0691_ _3276_ net124 sky130_fd_sc_hd__a32o_1
XFILLER_0_49_647 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6875_ VPWR VGND VPWR VGND _0465_ _2066_ _3242_ _3239_ _3051_ sky130_fd_sc_hd__a211oi_1
X_5826_ VGND VPWR VGND VPWR _2452_ _2088_ _2434_ net69 net81 sky130_fd_sc_hd__a211o_1
X_5757_ VPWR VGND VGND VPWR _2399_ _2398_ _2396_ sky130_fd_sc_hd__nor2_4
X_8545_ i_tinyqv.cpu.i_core.i_cycles.register\[18\] clknet_leaf_5_clk i_tinyqv.cpu.i_core.i_cycles.reg_buf\[18\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4708_ VPWR VGND VPWR VGND _1544_ net6 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_62_Left_143 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_8476_ VGND VPWR VGND VPWR i_tinyqv.cpu.debug_instr_valid _0574_ clknet_leaf_23_clk
+ sky130_fd_sc_hd__dfxtp_4
X_5688_ VGND VPWR VGND VPWR _0175_ net98 _2330_ _2346_ _2299_ sky130_fd_sc_hd__o211a_1
X_7427_ VPWR VGND _3675_ _3661_ i_tinyqv.cpu.instr_data_start\[11\] _0726_ i_tinyqv.cpu.instr_data_start\[13\]
+ VGND VPWR sky130_fd_sc_hd__a31o_1
X_4639_ VGND VPWR VPWR VGND _1475_ i_tinyqv.cpu.instr_data\[2\]\[14\] net322 i_tinyqv.cpu.instr_data\[0\]\[14\]
+ sky130_fd_sc_hd__mux2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.i_regbuf\[28\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[28\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_471 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_20_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7358_ VPWR VGND VGND VPWR _1405_ _3618_ _2147_ sky130_fd_sc_hd__nand2_1
X_6309_ VGND VPWR VPWR VGND _2765_ _2320_ _2762_ net269 sky130_fd_sc_hd__mux2_1
X_7289_ VPWR VGND VPWR VGND _3564_ _3563_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_71_Left_152 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_39_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_80_Left_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_23_536 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_4_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4990_ VPWR VGND VPWR VGND _1754_ i_tinyqv.cpu.no_write_in_progress sky130_fd_sc_hd__inv_2
X_3941_ VGND VPWR VPWR VGND _0792_ _0791_ _0790_ _0789_ _0793_ sky130_fd_sc_hd__or4_4
X_6660_ VGND VPWR VGND VPWR _3048_ _3040_ _3045_ _3046_ _3047_ sky130_fd_sc_hd__o211a_1
X_3872_ VPWR VGND VGND VPWR _0608_ _0724_ _0614_ sky130_fd_sc_hd__nand2_4
X_5611_ VPWR VGND VPWR VGND _2292_ _2281_ sky130_fd_sc_hd__inv_2
X_6591_ VPWR VGND _2989_ i_tinyqv.cpu.is_branch _0653_ VPWR VGND sky130_fd_sc_hd__and2_1
X_5542_ VGND VPWR net307 _2242_ _2244_ net91 VPWR VGND sky130_fd_sc_hd__o21ai_1
X_8330_ i_tinyqv.cpu.instr_fetch_stopped clknet_leaf_17_clk _0429_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5473_ VGND VPWR VPWR VGND _2193_ i_uart_tx.data_to_send\[7\] _2177_ i_uart_tx.data_to_send\[6\]
+ sky130_fd_sc_hd__mux2_1
X_8261_ i_tinyqv.cpu.instr_data_in\[1\] clknet_leaf_13_clk _0360_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_7212_ VGND VPWR VGND VPWR _3506_ i_tinyqv.cpu.instr_data\[2\]\[3\] _1432_ _1445_
+ _3489_ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_8192_ i_tinyqv.cpu.i_core.i_shift.a\[11\] clknet_leaf_41_clk _0304_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
X_4424_ VGND VPWR VPWR VGND _1267_ _1063_ _1088_ _1115_ sky130_fd_sc_hd__mux2_1
X_4355_ VPWR VGND VPWR VGND i_tinyqv.cpu.i_core.mcause\[1\] _0947_ _1198_ _0929_ i_tinyqv.cpu.i_core.i_instrret.data\[1\]
+ _1197_ sky130_fd_sc_hd__a221o_1
X_7143_ VGND VPWR VPWR VGND _3446_ _3447_ _3445_ _3448_ sky130_fd_sc_hd__or3b_1
X_7074_ VPWR VGND VPWR VGND _3385_ _2140_ _3382_ _3386_ _3364_ sky130_fd_sc_hd__a22o_1
X_4286_ VPWR VGND VGND VPWR _1080_ _1133_ _1132_ sky130_fd_sc_hd__nand2_1
X_6025_ VGND VPWR _0279_ _2578_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7976_ i_uart_tx.data_to_send\[3\] clknet_leaf_28_clk _0111_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_230 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_6927_ VGND VPWR VPWR VGND _0488_ _3269_ _3264_ _1589_ _3271_ net125 sky130_fd_sc_hd__a32o_1
X_6858_ VGND VPWR VPWR VGND _3224_ _3228_ _3227_ sky130_fd_sc_hd__xor2_1
X_5809_ VPWR VGND VPWR VGND _2438_ i_tinyqv.cpu.i_core.last_interrupt_req\[1\] sky130_fd_sc_hd__inv_2
XFILLER_0_9_574 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_29_190 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_6789_ _3165_ _3155_ _3147_ _3156_ _3153_ VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_8528_ i_tinyqv.cpu.i_core.i_cycles.register\[2\] clknet_leaf_4_clk _0598_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.i_regbuf\[29\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[29\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[1\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_8459_ i_tinyqv.cpu.i_core.mem_op\[1\] clknet_leaf_8_clk _0557_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_27_149 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_51_642 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.i_regbuf\[28\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[28\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_50_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_cycles.i_regbuf\[26\] i_tinyqv.cpu.i_core.i_cycles.reg_buf\[26\]
+ i_tinyqv.cpu.i_core.i_cycles.register\[30\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4140_ VPWR VGND _0987_ _0967_ i_tinyqv.cpu.data_addr\[4\] VPWR VGND sky130_fd_sc_hd__and2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.i_regbuf\[17\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[17\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[21\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4071_ VPWR VGND VPWR VGND _0917_ _0903_ _0858_ _0918_ sky130_fd_sc_hd__a21o_1
X_7830_ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[17\] clknet_leaf_3_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[17\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4973_ VGND VPWR _1744_ gpio_out_sel\[1\] _1737_ _1742_ VPWR VGND sky130_fd_sc_hd__and3_1
X_7761_ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[12\] clknet_leaf_1_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[12\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6712_ VGND VPWR VPWR VGND _3084_ _3087_ _3095_ _3085_ sky130_fd_sc_hd__a21boi_2
X_3924_ VPWR VGND VPWR VGND i_tinyqv.cpu.i_core.imm_lo\[5\] _0748_ _0776_ _0690_ i_tinyqv.cpu.i_core.imm_lo\[9\]
+ _0775_ sky130_fd_sc_hd__a221o_1
X_7692_ i_tinyqv.cpu.i_core.i_registers.reg_access\[10\]\[3\] clknet_leaf_57_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[7\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6643_ VGND VPWR _0443_ _3032_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_3855_ VGND VPWR VGND VPWR _0704_ _0703_ _0706_ _0707_ sky130_fd_sc_hd__o21bai_4
X_6574_ VPWR VGND VGND VPWR _2979_ i_tinyqv.mem.q_ctrl.spi_ram_a_select _2229_ sky130_fd_sc_hd__or2_1
X_3786_ VGND VPWR VGND VPWR _0627_ _0625_ _0626_ _0638_ _0624_ sky130_fd_sc_hd__nor4b_2
X_8313_ i_tinyqv.mem.q_ctrl.spi_in_buffer\[1\] clknet_leaf_15_clk _0412_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5525_ VGND VPWR _2230_ i_uart_tx.fsm_state\[0\] i_uart_tx.fsm_state\[1\] _2175_
+ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_74_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5456_ VGND VPWR _2181_ _2182_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_8244_ i_tinyqv.cpu.i_core.mepc\[15\] clknet_leaf_35_clk _0344_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_4407_ VPWR VGND VGND VPWR net68 _1250_ _0842_ sky130_fd_sc_hd__nor2_2
XFILLER_0_10_561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5387_ VGND VPWR _0103_ _2117_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8175_ i_tinyqv.cpu.instr_data\[1\]\[10\] clknet_leaf_10_clk _0287_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_4338_ VGND VPWR _1184_ i_tinyqv.cpu.debug_rd\[0\] VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_7126_ VGND VPWR _0526_ _3432_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4269_ VGND VPWR VPWR VGND _1116_ _1115_ _1108_ _1112_ sky130_fd_sc_hd__mux2_1
X_7057_ VGND VPWR _1461_ _3370_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_6008_ VGND VPWR VPWR VGND _2570_ i_tinyqv.cpu.instr_data\[2\]\[8\] _2563_ _2316_
+ sky130_fd_sc_hd__mux2_1
X_7959_ i_tinyqv.cpu.i_core.last_interrupt_req\[1\] clknet_leaf_26_clk _0096_ VPWR
+ VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_414 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_32_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_6290_ VGND VPWR _0368_ _2754_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_483 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5310_ VPWR VGND VGND VPWR _2057_ _0744_ _2056_ sky130_fd_sc_hd__nand2_2
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.i_regbuf\[18\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[18\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[22\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5241_ VPWR VGND _1995_ _1994_ _1993_ VPWR VGND sky130_fd_sc_hd__and2_1
X_5172_ VGND VPWR VPWR VGND _1926_ _1928_ _1927_ sky130_fd_sc_hd__xor2_1
X_4123_ _0970_ _0967_ i_tinyqv.cpu.data_addr\[4\] VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
Xinput2 VGND VPWR net2 ui_in[0] VPWR VGND sky130_fd_sc_hd__buf_1
X_4054_ VPWR VGND VGND VPWR i_tinyqv.cpu.instr_data_start\[20\] _0899_ _0901_ sky130_fd_sc_hd__nor2_1
X_7813_ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[0\] clknet_leaf_5_clk _0070_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_561 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7744_ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[27\] clknet_leaf_54_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[27\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_4956_ VPWR VGND VPWR VGND _1727_ net98 _1733_ _0002_ sky130_fd_sc_hd__a21o_1
X_7675_ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[22\] clknet_leaf_58_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[22\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.i_regbuf\[21\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[21\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[25\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3907_ VPWR VGND VPWR VGND _0637_ i_tinyqv.cpu.i_core.i_registers.reg_access\[7\]\[1\]
+ net88 _0759_ i_tinyqv.cpu.i_core.i_registers.reg_access\[11\]\[1\] sky130_fd_sc_hd__a22o_1
X_4887_ VGND VPWR VPWR VGND _1687_ _1303_ _1685_ i_tinyqv.cpu.i_core.i_registers.reg_access\[6\]\[1\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6626_ VPWR VGND VGND VPWR i_tinyqv.cpu.instr_data_start\[3\] _3019_ i_tinyqv.cpu.i_core.imm_lo\[3\]
+ sky130_fd_sc_hd__nand2_1
X_3838_ VGND VPWR _0620_ _0690_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_288 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_6557_ VGND VPWR _0424_ _2965_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5508_ VGND VPWR _0124_ _2217_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_3769_ VPWR VGND VPWR VGND _0620_ i_tinyqv.cpu.instr_data_start\[7\] _0619_ _0621_
+ i_tinyqv.cpu.instr_data_start\[11\] sky130_fd_sc_hd__a22o_1
X_6488_ VGND VPWR VPWR VGND _2904_ net271 _2897_ i_tinyqv.mem.q_ctrl.spi_in_buffer\[2\]
+ sky130_fd_sc_hd__mux2_1
X_8227_ i_tinyqv.cpu.i_core.multiplier.accum\[10\] clknet_leaf_43_clk _0017_ VPWR
+ VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.i_regbuf\[10\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[10\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[14\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5439_ _2166_ _2134_ _2136_ _2143_ _2165_ VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_8158_ i_tinyqv.cpu.instr_data\[2\]\[7\] clknet_leaf_10_clk _0270_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_7109_ VPWR VGND VPWR VGND i_tinyqv.cpu.instr_data\[3\]\[9\] _3369_ _3417_ _3370_
+ i_tinyqv.cpu.instr_data\[2\]\[9\] _3372_ sky130_fd_sc_hd__a221o_1
X_8089_ gpio_out\[0\] clknet_leaf_27_clk _0000_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_299 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_80_589 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_20_177 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4810_ VGND VPWR VPWR VGND _1643_ i_tinyqv.cpu.debug_rd\[0\] _1642_ i_tinyqv.cpu.i_core.i_registers.reg_access\[14\]\[0\]
+ sky130_fd_sc_hd__mux2_1
X_5790_ VPWR VGND _2424_ _2423_ _2181_ VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_8_628 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_4741_ VGND VPWR _1576_ _1315_ _1575_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_22_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_71_512 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7460_ VGND VPWR VPWR VGND _3703_ _3702_ _3239_ _3190_ sky130_fd_sc_hd__mux2_1
X_4672_ VGND VPWR VPWR VGND _1508_ i_tinyqv.cpu.instr_data\[3\]\[7\] _1449_ i_tinyqv.cpu.instr_data\[1\]\[7\]
+ sky130_fd_sc_hd__mux2_1
X_6411_ _2847_ _1706_ _2846_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_7391_ VGND VPWR _3645_ _0883_ i_tinyqv.cpu.instr_data_start\[7\] _3634_ VPWR VGND
+ sky130_fd_sc_hd__and3_1
X_6342_ VPWR VGND VGND VPWR i_tinyqv.mem.data_stall _1532_ _2783_ sky130_fd_sc_hd__or2b_2
X_6273_ VGND VPWR VPWR VGND _2746_ i_tinyqv.cpu.instr_data_in\[1\] _2744_ _2318_ sky130_fd_sc_hd__mux2_1
X_8012_ i_uart_rx.recieved_data\[5\] clknet_leaf_19_clk _0147_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_5224_ VGND VPWR VPWR VGND _1976_ _1978_ _1977_ sky130_fd_sc_hd__xor2_1
X_5155_ VPWR VGND VGND VPWR _1910_ _1912_ _1911_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5086_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[6\] _1846_ _1845_ sky130_fd_sc_hd__nand2_1
X_4106_ VPWR VGND VPWR VGND _0918_ _0707_ _0880_ _0953_ _0952_ sky130_fd_sc_hd__a22o_1
X_4037_ VPWR VGND _0884_ i_tinyqv.cpu.instr_data_start\[3\] VPWR VGND sky130_fd_sc_hd__buf_2
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.i_regbuf\[22\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[22\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[26\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5988_ VPWR VGND _2558_ _2557_ _2079_ VPWR VGND sky130_fd_sc_hd__and2_1
X_4939_ VPWR VGND _1721_ i_tinyqv.cpu.instr_data_in\[15\] VPWR VGND sky130_fd_sc_hd__buf_2
X_7727_ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[10\] clknet_leaf_0_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[10\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XANTENNA_40 i_tinyqv.cpu.i_core.imm_lo\[9\] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_7658_ i_tinyqv.cpu.i_core.i_registers.reg_access\[11\]\[1\] clknet_leaf_55_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[5\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6609_ VGND VPWR _3004_ _3005_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.i_regbuf\[8\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[8\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[12\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_62_589 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7589_ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[0\] clknet_leaf_57_clk _0046_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.i_regbuf\[11\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[11\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[15\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.i_regbuf\[18\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[18\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[22\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.i_regbuf\[6\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[6\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[10\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_72_309 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_25_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_53_545 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_4_108 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_80_386 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.i_regbuf\[10\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[10\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[14\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6960_ VPWR VGND VPWR VGND _1483_ _1487_ _1468_ _3283_ sky130_fd_sc_hd__or3_1
X_5911_ VGND VPWR VPWR VGND _2506_ _2505_ _2502_ net137 sky130_fd_sc_hd__mux2_1
XFILLER_0_17_96 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6891_ VPWR VGND _0471_ _3251_ _3243_ _1387_ _3252_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_5842_ VPWR VGND _2463_ _2462_ VPWR VGND sky130_fd_sc_hd__buf_4
X_5773_ VPWR VGND VPWR VGND _2411_ i_spi.bits_remaining\[2\] _2406_ _2412_ _2404_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_414 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_8561_ i_tinyqv.cpu.i_core.i_instrret.register\[0\] clknet_leaf_50_clk _0603_ VPWR
+ VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_73 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_33_95 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_4724_ VGND VPWR _1559_ net8 _1560_ net7 VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_7512_ VGND VPWR _3745_ i_tinyqv.cpu.i_core.i_instrret.data\[1\] net92 _3744_ VPWR
+ VGND sky130_fd_sc_hd__and3_1
XFILLER_0_71_331 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_8492_ i_tinyqv.mem.q_ctrl.addr\[18\] clknet_leaf_32_clk _0590_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_7443_ VGND VPWR VGND VPWR _3689_ net173 _3012_ _3004_ _3688_ sky130_fd_sc_hd__o211a_1
X_4655_ VGND VPWR VGND VPWR _1462_ _1416_ _1464_ _1491_ sky130_fd_sc_hd__a21o_2
X_7374_ VPWR VGND VGND VPWR net310 _3624_ _2733_ _3631_ sky130_fd_sc_hd__o21a_1
X_4586_ VPWR VGND _1422_ _1417_ VPWR VGND sky130_fd_sc_hd__buf_2
X_6325_ VGND VPWR VPWR VGND _2774_ _2318_ _2772_ net286 sky130_fd_sc_hd__mux2_1
XFILLER_0_4_697 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6256_ VGND VPWR VGND VPWR _2732_ _1541_ _1551_ _1536_ sky130_fd_sc_hd__a21o_4
X_5207_ VPWR VGND VGND VPWR _1960_ _1962_ _1961_ sky130_fd_sc_hd__nand2_1
X_6187_ VGND VPWR _0345_ _2674_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5138_ VGND VPWR _1867_ _1895_ _1896_ _1866_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_5069_ VPWR VGND VGND VPWR _1827_ _1829_ _0020_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_30_283 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_38_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_58_604 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.i_regbuf\[22\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[22\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[26\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_38_394 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_26_589 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xhold107 net136 i_tinyqv.cpu.data_out\[13\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4440_ VGND VPWR VPWR VGND _1283_ _1138_ _1108_ _1135_ sky130_fd_sc_hd__mux2_1
Xhold118 net147 i_tinyqv.mem.q_ctrl.addr\[12\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 net158 i_tinyqv.cpu.i_core.mcause\[4\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6110_ VGND VPWR VPWR VGND _2623_ i_tinyqv.cpu.i_core.i_shift.a\[27\] _2595_ i_tinyqv.cpu.i_core.i_shift.a\[31\]
+ sky130_fd_sc_hd__mux2_1
X_4371_ VGND VPWR VPWR VGND _1214_ _0610_ _1211_ _0916_ _1213_ sky130_fd_sc_hd__o2bb2a_1
X_7090_ VPWR VGND VGND VPWR _3398_ _3399_ _3304_ _3400_ sky130_fd_sc_hd__o21a_1
X_6041_ VGND VPWR _0287_ _2586_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7992_ i_uart_tx.fsm_state\[0\] clknet_leaf_32_clk _0127_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_6943_ VGND VPWR VPWR VGND _0499_ _3274_ _3268_ _0691_ _3276_ net119 sky130_fd_sc_hd__a32o_1
X_6874_ VGND VPWR VGND VPWR _3051_ _1550_ _3241_ _3242_ sky130_fd_sc_hd__o21ba_1
X_5825_ VPWR VGND VGND VPWR net179 _2451_ _2450_ sky130_fd_sc_hd__nand2_1
X_5756_ VPWR VGND VGND VPWR i_spi.spi_clk_out _2384_ _2398_ sky130_fd_sc_hd__nor2_1
X_8544_ i_tinyqv.cpu.i_core.i_cycles.register\[17\] clknet_leaf_4_clk i_tinyqv.cpu.i_core.i_cycles.reg_buf\[17\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5687_ VGND VPWR VGND VPWR _2346_ _2336_ _2341_ net255 _2345_ sky130_fd_sc_hd__a211o_1
X_4707_ VGND VPWR VGND VPWR _1543_ _1542_ _1534_ i_tinyqv.mem.instr_active _1537_
+ sky130_fd_sc_hd__a31o_4
X_8475_ i_tinyqv.cpu.i_core.is_interrupt clknet_leaf_7_clk _0573_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_2
X_7426_ VPWR VGND VGND VPWR _3625_ net147 _3624_ net153 _0584_ _3674_ sky130_fd_sc_hd__o221a_1
X_4638_ VGND VPWR VPWR VGND _1474_ i_tinyqv.cpu.instr_data\[3\]\[14\] net322 i_tinyqv.cpu.instr_data\[1\]\[14\]
+ sky130_fd_sc_hd__mux2_1
X_7357_ VPWR VGND VGND VPWR _3312_ _3474_ i_tinyqv.cpu.mem_op_increment_reg _3617_
+ _0572_ sky130_fd_sc_hd__o22a_1
X_4569_ VPWR VGND VGND VPWR _0862_ _1404_ _1405_ sky130_fd_sc_hd__nor2_1
X_6308_ VGND VPWR _0376_ _2764_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7288_ VPWR VGND VPWR VGND _3553_ _3299_ _3562_ _3563_ sky130_fd_sc_hd__a21o_1
X_6239_ VGND VPWR VPWR VGND _2716_ _2718_ _2717_ sky130_fd_sc_hd__xor2_1
X_3940_ VPWR VGND VPWR VGND net48 i_tinyqv.cpu.i_core.i_registers.reg_access\[1\]\[2\]
+ _0648_ _0792_ i_tinyqv.cpu.i_core.i_registers.reg_access\[14\]\[2\] sky130_fd_sc_hd__a22o_1
X_3871_ VGND VPWR _0723_ _0611_ i_tinyqv.cpu.instr_data_start\[8\] _0690_ VPWR VGND
+ sky130_fd_sc_hd__and3_1
X_5610_ VPWR VGND VPWR VGND _2285_ _1228_ _2282_ _2291_ _2278_ sky130_fd_sc_hd__a22o_1
X_6590_ VGND VPWR VPWR VGND _0749_ _2988_ i_tinyqv.cpu.i_core.imm_lo\[1\] sky130_fd_sc_hd__xor2_1
XFILLER_0_6_704 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_5541_ VGND VPWR _0131_ _2243_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_651 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_5_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_8260_ i_tinyqv.cpu.instr_data_in\[0\] clknet_leaf_13_clk _0359_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_5472_ VGND VPWR VGND VPWR _0113_ i_debug_uart_tx.uart_tx_data\[5\] _2169_ _2192_
+ _2182_ sky130_fd_sc_hd__o211a_1
X_7211_ VPWR VGND VGND VPWR i_tinyqv.cpu.imm\[18\] _3360_ _3505_ _0538_ sky130_fd_sc_hd__o21a_1
XFILLER_0_10_710 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_8191_ i_tinyqv.cpu.i_core.i_shift.a\[10\] clknet_leaf_41_clk _0303_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
X_4423_ VGND VPWR VPWR VGND _1266_ _1112_ _1149_ _1107_ sky130_fd_sc_hd__mux2_1
X_4354_ VPWR VGND VPWR VGND _1196_ i_tinyqv.cpu.i_core.cycle_count\[1\] _0931_ _1197_
+ _0927_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_50 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_7142_ VGND VPWR _3337_ _3298_ _3447_ _2130_ VPWR VGND sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_18_Left_99 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7073_ VGND VPWR VPWR VGND _3385_ _3384_ _3319_ _1514_ sky130_fd_sc_hd__mux2_1
X_6024_ VGND VPWR VPWR VGND _2578_ i_tinyqv.cpu.instr_data\[1\]\[2\] _2463_ i_tinyqv.cpu.instr_data_in\[2\]
+ sky130_fd_sc_hd__mux2_1
X_4285_ VGND VPWR VPWR VGND _1132_ _1131_ _1088_ _1130_ sky130_fd_sc_hd__mux2_1
X_7975_ i_uart_tx.data_to_send\[2\] clknet_leaf_29_clk _0110_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_6926_ VGND VPWR VPWR VGND _0487_ _3268_ _3264_ _1589_ _3271_ net130 sky130_fd_sc_hd__a32o_1
X_6857_ VGND VPWR VGND VPWR _3225_ _3227_ _3226_ sky130_fd_sc_hd__or2b_1
X_6788_ VPWR VGND VPWR VGND _3164_ net105 sky130_fd_sc_hd__inv_2
X_5808_ VGND VPWR _2102_ _0613_ _2437_ net66 VPWR VGND sky130_fd_sc_hd__o21ai_1
X_5739_ VPWR VGND VPWR VGND _2381_ _2380_ _2382_ _2383_ sky130_fd_sc_hd__a21oi_1
X_8527_ i_tinyqv.cpu.i_core.i_cycles.register\[1\] clknet_leaf_3_clk _0597_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_8458_ VGND VPWR VGND VPWR i_tinyqv.cpu.i_core.mem_op\[0\] _0556_ clknet_leaf_6_clk
+ sky130_fd_sc_hd__dfxtp_4
X_8389_ i_tinyqv.cpu.data_out\[14\] clknet_leaf_19_clk _0487_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_7409_ VPWR VGND VGND VPWR _3239_ _3108_ _3660_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_570 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.i_regbuf\[25\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[25\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[29\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_cycles.i_regbuf\[19\] i_tinyqv.cpu.i_core.i_cycles.reg_buf\[19\]
+ i_tinyqv.cpu.i_core.i_cycles.register\[23\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4070_ VPWR VGND VGND VPWR _0916_ _0913_ _0688_ _0915_ _0917_ sky130_fd_sc_hd__o22a_1
X_4972_ VPWR VGND VPWR VGND _1741_ net117 _1743_ _0008_ sky130_fd_sc_hd__a21o_1
X_7760_ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[11\] clknet_leaf_57_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[11\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6711_ VGND VPWR VPWR VGND _3094_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[17\]
+ net31 _1202_ sky130_fd_sc_hd__mux2_1
X_3923_ VGND VPWR _0775_ _0608_ _0614_ i_tinyqv.cpu.imm\[13\] VPWR VGND sky130_fd_sc_hd__and3_1
X_7691_ i_tinyqv.cpu.i_core.i_registers.reg_access\[10\]\[2\] clknet_leaf_53_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[6\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_212 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_6642_ VGND VPWR VPWR VGND _3032_ net308 _2415_ i_spi.end_txn sky130_fd_sc_hd__mux2_1
X_3854_ VPWR VGND VGND VPWR _0611_ _0705_ _0706_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_673 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_8312_ i_tinyqv.mem.q_ctrl.spi_in_buffer\[0\] clknet_leaf_16_clk _0411_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6573_ VGND VPWR _0427_ _2978_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_3785_ VPWR VGND VGND VPWR _0625_ net324 _0627_ _0624_ _0637_ sky130_fd_sc_hd__and4b_2
X_5524_ VGND VPWR _2198_ _2229_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_5455_ VGND VPWR _1728_ _2181_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_8243_ i_tinyqv.cpu.i_core.mepc\[14\] clknet_leaf_34_clk _0343_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_4406_ VPWR VGND VGND VPWR _1247_ _1249_ _1248_ sky130_fd_sc_hd__nand2_1
X_8174_ i_tinyqv.cpu.instr_data\[1\]\[9\] clknet_leaf_10_clk _0286_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5386_ VPWR VGND VGND VPWR _2117_ _2083_ _2116_ sky130_fd_sc_hd__or2_1
X_7125_ VGND VPWR VPWR VGND _3432_ _3431_ _3396_ i_tinyqv.cpu.i_core.imm_lo\[6\] sky130_fd_sc_hd__mux2_1
X_4337_ VGND VPWR VPWR VGND _1184_ _1024_ _0954_ _0877_ _1035_ _1183_ sky130_fd_sc_hd__a32o_1
X_4268_ VGND VPWR VPWR VGND _1115_ _1114_ _1050_ _1113_ sky130_fd_sc_hd__mux2_1
X_7056_ VGND VPWR _1504_ _3369_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_6007_ VGND VPWR _0270_ _2569_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4199_ VGND VPWR VPWR VGND _1045_ _1044_ _1046_ _1038_ sky130_fd_sc_hd__a21boi_2
X_7958_ i_tinyqv.cpu.i_core.last_interrupt_req\[0\] clknet_leaf_26_clk _0095_ VPWR
+ VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6909_ VPWR VGND _3265_ _3264_ VPWR VGND sky130_fd_sc_hd__buf_2
X_7889_ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[12\] clknet_leaf_49_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[12\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_275 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_37_437 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xhold290 net319 i_debug_uart_tx.uart_tx_data\[6\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.i_regbuf\[26\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[26\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[30\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_43_429 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_11_326 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_5240_ VPWR VGND VGND VPWR _1994_ _1991_ _1992_ sky130_fd_sc_hd__or2_1
X_5171_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[11\] _1927_ _1167_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_18_Right_18 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4122_ VPWR VGND VPWR VGND _0961_ _0966_ i_tinyqv.cpu.data_addr\[3\] _0969_ sky130_fd_sc_hd__or3_4
X_4053_ VPWR VGND _0900_ _0899_ i_tinyqv.cpu.instr_data_start\[20\] VPWR VGND sky130_fd_sc_hd__and2_1
Xinput3 VGND VPWR net3 ui_in[1] VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7812_ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[31\] clknet_leaf_0_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[31\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4955_ VGND VPWR _1733_ gpio_out\[2\] _1729_ _1730_ VPWR VGND sky130_fd_sc_hd__and3_1
X_7743_ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[26\] clknet_leaf_0_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[26\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_404 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_27_Right_27 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_74_510 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_3906_ VPWR VGND VPWR VGND _0639_ i_tinyqv.cpu.i_core.i_registers.reg_access\[5\]\[1\]
+ net57 _0758_ i_tinyqv.cpu.i_core.i_registers.reg_access\[6\]\[1\] sky130_fd_sc_hd__a22o_1
X_7674_ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[21\] clknet_leaf_55_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[21\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4886_ VGND VPWR _0066_ _1686_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6625_ VPWR VGND VPWR VGND i_tinyqv.cpu.instr_write_offset\[3\] _0884_ _3017_ _3018_
+ sky130_fd_sc_hd__a21oi_1
X_3837_ VPWR VGND _0689_ _0615_ VPWR VGND sky130_fd_sc_hd__buf_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.i_regbuf\[14\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[14\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[18\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6556_ VGND VPWR VPWR VGND _2965_ _1717_ _2925_ _2964_ sky130_fd_sc_hd__mux2_1
X_3768_ VGND VPWR VPWR VGND i_tinyqv.cpu.counter\[2\] _0620_ i_tinyqv.cpu.counter\[3\]
+ sky130_fd_sc_hd__and2b_2
XFILLER_0_15_643 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5507_ _2215_ _2199_ _2217_ _2216_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_6487_ VGND VPWR _0416_ net134 VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8226_ i_tinyqv.cpu.i_core.multiplier.accum\[9\] clknet_leaf_44_clk _0027_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_36_Right_36 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5438_ VGND VPWR _1498_ _2165_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_8157_ i_tinyqv.cpu.instr_data\[2\]\[6\] clknet_leaf_4_clk _0269_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5369_ VPWR VGND VPWR VGND net69 _0656_ _1185_ _2102_ sky130_fd_sc_hd__a21o_1
X_8088_ gpio_out_sel\[7\] clknet_leaf_17_clk _0015_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7108_ VPWR VGND VGND VPWR _3347_ _3416_ _3415_ sky130_fd_sc_hd__nand2_1
X_7039_ VPWR VGND VGND VPWR _3353_ _3292_ _3284_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_45_Right_45 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_54_Right_54 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_63_Right_63 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4740_ VPWR VGND _1575_ _1574_ _1573_ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_28_234 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.i_regbuf\[9\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[9\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[13\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4671_ VGND VPWR VGND VPWR _1503_ _1506_ _1507_ _1461_ sky130_fd_sc_hd__a21oi_4
X_6410_ VPWR VGND _2846_ _1707_ i_tinyqv.mem.q_ctrl.fsm_state\[1\] VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_71_557 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7390_ VPWR VGND VGND VPWR _3644_ _3625_ net89 _3643_ _0578_ sky130_fd_sc_hd__o22a_1
XFILLER_0_43_248 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6341_ VPWR VGND VGND VPWR _2782_ i_tinyqv.mem.q_ctrl.read_cycles_count\[1\] i_tinyqv.mem.q_ctrl.read_cycles_count\[2\]
+ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_72_Right_72 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_12_602 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.i_regbuf\[30\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[30\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[2\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6272_ VGND VPWR _0359_ _2745_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8011_ i_uart_rx.recieved_data\[4\] clknet_leaf_18_clk _0146_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_5223_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[13\] _1977_ _1167_ sky130_fd_sc_hd__nand2_1
X_5154_ VPWR VGND VGND VPWR _1911_ i_tinyqv.cpu.i_core.multiplier.accum\[10\] _1909_
+ sky130_fd_sc_hd__or2_1
X_4105_ VPWR VGND VPWR VGND _0951_ _0921_ _0880_ _0952_ sky130_fd_sc_hd__a21oi_1
X_5085_ VGND VPWR _1250_ _1845_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_613 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4036_ VPWR VGND _0883_ i_tinyqv.cpu.instr_data_start\[6\] VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_0_2_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5987_ VPWR VGND VPWR VGND _2552_ i_tinyqv.cpu.data_addr\[26\] _1758_ _2557_ i_tinyqv.cpu.i_core.i_shift.a\[30\]
+ sky130_fd_sc_hd__a22o_1
X_4938_ VGND VPWR VGND VPWR uio_out[4] _1720_ i_tinyqv.mem.q_ctrl.addr\[22\] _1709_
+ _1711_ sky130_fd_sc_hd__a22o_4
X_7726_ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[9\] clknet_leaf_54_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[9\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.i_regbuf\[15\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[15\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[19\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_30 i_tinyqv.cpu.i_core.imm_lo\[4\] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_41 i_tinyqv.cpu.i_core.imm_lo\[9\] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_7657_ i_tinyqv.cpu.i_core.i_registers.reg_access\[11\]\[0\] clknet_leaf_1_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[4\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4869_ VGND VPWR _0075_ _1676_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6608_ VGND VPWR VGND VPWR _1536_ _1541_ _3004_ _1551_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_62_557 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_7588_ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[31\] clknet_leaf_59_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[31\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6539_ VGND VPWR VPWR VGND _2950_ _2949_ _2792_ _2947_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_30_432 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_8209_ i_tinyqv.cpu.i_core.i_shift.a\[30\] clknet_leaf_39_clk _0321_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.i_regbuf\[8\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[8\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[12\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap21 VGND VPWR net21 net22 VPWR VGND sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_6_Left_87 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_43_19 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_80_365 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.i_regbuf\[6\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[6\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[10\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5910_ VGND VPWR VPWR VGND _2504_ i_tinyqv.cpu.i_core.mepc\[1\] i_tinyqv.cpu.i_core.i_shift.a\[5\]
+ _2505_ sky130_fd_sc_hd__mux2_2
X_6890_ VPWR VGND VPWR VGND _1604_ i_tinyqv.cpu.no_write_in_progress _2066_ _3252_
+ sky130_fd_sc_hd__a21o_1
X_5841_ VGND VPWR _2461_ _2462_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_5772_ VGND VPWR _2402_ _2411_ i_spi.bits_remaining\[2\] VPWR VGND sky130_fd_sc_hd__xnor2_1
X_8560_ i_tinyqv.cpu.i_core.i_cycles.cy clknet_leaf_51_clk _0602_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_8491_ i_tinyqv.mem.q_ctrl.addr\[17\] clknet_leaf_32_clk _0589_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_4723_ VGND VPWR VGND VPWR _1556_ _1555_ net5 _1558_ _1557_ net6 _1559_ sky130_fd_sc_hd__mux4_1
X_7511_ VGND VPWR VPWR VGND _3744_ i_tinyqv.cpu.i_core.i_instrret.cy _1026_ i_tinyqv.cpu.i_core.i_instrret.add
+ sky130_fd_sc_hd__mux2_1
X_7442_ VPWR VGND VPWR VGND _3632_ _3158_ _3688_ _3686_ _3687_ _2877_ sky130_fd_sc_hd__a221o_1
XFILLER_0_71_354 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4654_ VGND VPWR _1489_ _1490_ VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_0_44_568 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7373_ VPWR VGND VGND VPWR _3628_ _3629_ _3630_ sky130_fd_sc_hd__nor2_1
X_4585_ VPWR VGND VGND VPWR _1421_ i_tinyqv.cpu.instr_data\[1\]\[1\] _1414_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_218 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_6324_ VGND VPWR _0383_ _2773_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6255_ VPWR VGND _0356_ _2730_ _1813_ _1060_ _2731_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_5206_ VPWR VGND VGND VPWR _1961_ i_tinyqv.cpu.i_core.multiplier.accum\[12\] _1959_
+ sky130_fd_sc_hd__or2_1
X_6186_ VGND VPWR VPWR VGND _2674_ i_tinyqv.cpu.i_core.mepc\[20\] _2667_ i_tinyqv.cpu.i_core.mepc\[16\]
+ sky130_fd_sc_hd__mux2_1
X_5137_ VGND VPWR VGND VPWR _1864_ _1895_ _1865_ sky130_fd_sc_hd__or2b_1
X_5068_ VPWR VGND VGND VPWR _1825_ _1828_ _1829_ sky130_fd_sc_hd__nor2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.i_regbuf\[5\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[5\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[9\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4019_ VGND VPWR VGND VPWR i_tinyqv.cpu.data_write_n\[0\] i_tinyqv.cpu.data_read_n\[0\]
+ _0869_ _0866_ sky130_fd_sc_hd__a21oi_2
XPHY_EDGE_ROW_0_Right_0 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7709_ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[24\] clknet_leaf_2_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[24\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.i_regbuf\[30\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[30\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[2\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.i_regbuf\[15\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[15\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[19\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold108 net137 i_tinyqv.cpu.data_addr\[1\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold119 net148 i_uart_rx.cycle_counter\[4\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4370_ VPWR VGND VGND VPWR _1213_ _0898_ _1212_ sky130_fd_sc_hd__or2_1
X_6040_ VGND VPWR VPWR VGND _2586_ i_tinyqv.cpu.instr_data\[1\]\[10\] _2462_ _2320_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7991_ i_uart_tx.cycle_counter\[10\] clknet_leaf_31_clk _0126_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_6942_ VGND VPWR VPWR VGND _0498_ _3274_ _3267_ _0691_ _3276_ net118 sky130_fd_sc_hd__a32o_1
XFILLER_0_49_605 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6873_ VPWR VGND VPWR VGND _3240_ i_tinyqv.cpu.instr_fetch_running net183 _3241_
+ sky130_fd_sc_hd__a21oi_1
X_5824_ VPWR VGND VPWR VGND _2088_ net81 _2434_ _2450_ sky130_fd_sc_hd__a21o_1
X_5755_ VPWR VGND VGND VPWR i_spi.bits_remaining\[3\] _2396_ _2397_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_278 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_8543_ i_tinyqv.cpu.i_core.i_cycles.register\[16\] clknet_leaf_51_clk i_tinyqv.cpu.i_core.i_cycles.reg_buf\[16\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5686_ VPWR VGND _2345_ _2337_ i_debug_uart_tx.data_to_send\[3\] VPWR VGND sky130_fd_sc_hd__and2_1
X_4706_ VGND VPWR _1538_ _1541_ _1542_ i_tinyqv.mem.instr_active VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_568 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_8474_ i_tinyqv.cpu.mem_op_increment_reg clknet_leaf_6_clk _0572_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_7425_ VGND VPWR VGND VPWR _3674_ _2878_ _2732_ i_tinyqv.cpu.data_addr\[12\] _3673_
+ sky130_fd_sc_hd__a211o_1
X_4637_ VGND VPWR VGND VPWR _1470_ _1472_ _1473_ _1461_ sky130_fd_sc_hd__a21oi_4
X_7356_ VPWR VGND VGND VPWR _2079_ _3617_ _3562_ sky130_fd_sc_hd__nand2_1
X_4568_ VGND VPWR VGND VPWR _1404_ _1403_ _1402_ i_tinyqv.cpu.i_core.mstatus_mie sky130_fd_sc_hd__a21bo_1
X_6307_ VGND VPWR VPWR VGND _2764_ _2318_ _2762_ net277 sky130_fd_sc_hd__mux2_1
X_4499_ VPWR VGND VGND VPWR _0896_ _1337_ _1338_ sky130_fd_sc_hd__nor2_1
X_7287_ _3562_ _1507_ _2123_ _2124_ _3320_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
X_6238_ VGND VPWR _2717_ _1813_ i_tinyqv.cpu.i_core.i_shift.a\[14\] _2024_ VPWR VGND
+ sky130_fd_sc_hd__and3_1
X_6169_ VGND VPWR VPWR VGND _2665_ net228 _2656_ i_tinyqv.cpu.i_core.mepc\[8\] sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_20_clk VGND VPWR clknet_3_3__leaf_clk clknet_leaf_20_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_9_Left_90 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_3870_ VGND VPWR net77 _0658_ _0722_ _0708_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_5540_ _2243_ i_uart_rx.cycle_counter\[0\] _2242_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_11_clk VGND VPWR clknet_3_2__leaf_clk clknet_leaf_11_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_5471_ VPWR VGND VGND VPWR _2192_ _2179_ _2191_ sky130_fd_sc_hd__or2_1
X_4422_ VGND VPWR VGND VPWR _1265_ _1120_ _1092_ _1149_ _1264_ sky130_fd_sc_hd__a211o_1
X_7210_ VGND VPWR VGND VPWR _3505_ _3504_ _3500_ _3476_ _3438_ sky130_fd_sc_hd__a211o_1
X_8190_ i_tinyqv.cpu.i_core.i_shift.a\[9\] clknet_leaf_41_clk _0302_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
X_4353_ VGND VPWR VPWR VGND _1196_ i_tinyqv.cpu.i_core.cycle_count_wide\[4\] _0841_
+ i_tinyqv.cpu.i_core.time_hi\[0\] sky130_fd_sc_hd__mux2_1
X_7141_ VGND VPWR _3446_ _3299_ _2155_ _2120_ VPWR VGND sky130_fd_sc_hd__and3_1
X_4284_ VGND VPWR VPWR VGND _1131_ _1096_ _1083_ _1094_ sky130_fd_sc_hd__mux2_1
X_7072_ VPWR VGND VGND VPWR _3368_ i_tinyqv.cpu.instr_data\[1\]\[5\] _3366_ i_tinyqv.cpu.instr_data\[0\]\[5\]
+ _3384_ _3383_ sky130_fd_sc_hd__o221a_2
X_6023_ VGND VPWR _0278_ _2577_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7974_ i_uart_tx.data_to_send\[1\] clknet_leaf_29_clk _0109_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_6925_ VGND VPWR VPWR VGND _0486_ _3267_ _3265_ _1589_ _3271_ net136 sky130_fd_sc_hd__a32o_1
X_6856_ VPWR VGND VGND VPWR i_tinyqv.cpu.instr_data_start\[22\] _3226_ i_tinyqv.cpu.imm\[22\]
+ sky130_fd_sc_hd__nand2_1
X_6787_ VGND VPWR VGND VPWR _0456_ _0881_ _3123_ _3163_ _3093_ sky130_fd_sc_hd__o211a_1
X_3999_ VGND VPWR VGND VPWR _0850_ _0847_ _0849_ _0842_ i_tinyqv.cpu.i_core.cycle\[1\]
+ sky130_fd_sc_hd__a211o_1
X_5807_ VPWR VGND _2436_ _2088_ net66 _0613_ _2435_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_5738_ VGND VPWR VPWR VGND i_spi.clock_divider\[0\] _2382_ i_spi.clock_count\[0\]
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_17_332 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_8526_ i_tinyqv.cpu.i_core.i_cycles.register\[0\] clknet_leaf_6_clk _0596_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5669_ VPWR VGND _2330_ _2329_ VPWR VGND sky130_fd_sc_hd__buf_2
X_8457_ VGND VPWR VGND VPWR i_tinyqv.cpu.alu_op\[3\] _0555_ clknet_leaf_6_clk sky130_fd_sc_hd__dfxtp_4
X_8388_ i_tinyqv.cpu.data_out\[13\] clknet_leaf_19_clk _0486_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_7408_ VPWR VGND VPWR VGND net305 _3007_ _0581_ _3009_ net187 _3659_ sky130_fd_sc_hd__a221o_1
XFILLER_0_13_582 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_7339_ VGND VPWR _0566_ _3605_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.i_regbuf\[29\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[29\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[1\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.i_regbuf\[18\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[18\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[22\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xi_tinyqv.cpu.i_core.i_instrret.i_regbuf\[28\] i_tinyqv.cpu.i_core.i_instrret.reg_buf\[28\]
+ i_tinyqv.cpu.i_core.i_instrret.register\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_0_clk VGND VPWR clknet_3_0__leaf_clk clknet_leaf_0_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_4971_ VGND VPWR _1743_ gpio_out_sel\[0\] _1737_ _1742_ VPWR VGND sky130_fd_sc_hd__and3_1
X_6710_ VGND VPWR VGND VPWR _0449_ i_tinyqv.cpu.instr_data_start\[8\] _3027_ _3092_
+ _3093_ sky130_fd_sc_hd__o211a_1
X_7690_ i_tinyqv.cpu.i_core.i_registers.reg_access\[10\]\[1\] clknet_leaf_53_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[5\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_416 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_3922_ VPWR VGND VPWR VGND _0615_ i_tinyqv.cpu.i_core.imm_lo\[1\] i_tinyqv.cpu.counter\[4\]
+ _0774_ sky130_fd_sc_hd__a21o_1
X_6641_ VGND VPWR VGND VPWR _0442_ net60 _3027_ _3031_ _2061_ sky130_fd_sc_hd__o211a_1
X_3853_ VGND VPWR VGND VPWR i_tinyqv.cpu.imm\[20\] i_tinyqv.cpu.imm\[16\] _0608_ i_tinyqv.cpu.imm\[28\]
+ i_tinyqv.cpu.imm\[24\] _0614_ _0705_ sky130_fd_sc_hd__mux4_1
X_6572_ VPWR VGND VGND VPWR _2978_ net311 _2229_ sky130_fd_sc_hd__or2_1
X_3784_ VGND VPWR VGND VPWR net62 i_tinyqv.cpu.i_core.i_registers.reg_access\[13\]\[3\]
+ _0635_ _0636_ _0632_ sky130_fd_sc_hd__a211o_4
X_8311_ i_tinyqv.cpu.i_core.i_shift.a\[29\] clknet_leaf_39_clk _0410_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
X_5523_ VGND VPWR _0128_ _2228_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5454_ VPWR VGND VGND VPWR _2180_ _2178_ _2179_ sky130_fd_sc_hd__or2_1
X_8242_ i_tinyqv.cpu.i_core.mepc\[13\] clknet_leaf_35_clk _0342_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_4405_ VPWR VGND VGND VPWR _1169_ _1248_ _1246_ sky130_fd_sc_hd__nand2_1
X_5385_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.mstatus_mte _2107_ _2057_ _2116_ sky130_fd_sc_hd__o21a_1
X_8173_ i_tinyqv.cpu.instr_data\[1\]\[8\] clknet_leaf_11_clk _0285_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_4336_ VPWR VGND VPWR VGND _1033_ _1182_ _1165_ _1183_ sky130_fd_sc_hd__or3_1
X_7124_ VPWR VGND VPWR VGND _3425_ _3430_ _3429_ _3424_ _3431_ sky130_fd_sc_hd__or4_1
XFILLER_0_5_52 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4267_ VGND VPWR VPWR VGND _1114_ _1060_ _1036_ i_tinyqv.cpu.i_core.i_shift.a\[16\]
+ sky130_fd_sc_hd__mux2_1
X_7055_ VGND VPWR _3367_ _3368_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_4198_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.b\[4\] _1045_ _1037_ sky130_fd_sc_hd__nand2_1
X_6006_ VGND VPWR VPWR VGND _2569_ i_tinyqv.cpu.instr_data\[2\]\[7\] _2563_ i_tinyqv.cpu.instr_data_in\[7\]
+ sky130_fd_sc_hd__mux2_1
X_7957_ i_tinyqv.cpu.i_core.i_instrret.add clknet_leaf_50_clk net128 VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_6908_ VGND VPWR _3264_ i_tinyqv.cpu.no_write_in_progress i_tinyqv.cpu.is_store _3263_
+ VPWR VGND sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_59_Left_140 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7888_ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[11\] clknet_leaf_48_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[11\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_405 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_6839_ VGND VPWR VPWR VGND _3207_ _3211_ _3210_ sky130_fd_sc_hd__xor2_1
X_8509_ i_tinyqv.cpu.i_core.i_instrret.register\[15\] clknet_leaf_45_clk i_tinyqv.cpu.i_core.i_instrret.reg_buf\[15\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold280 net309 i_debug_uart_tx.uart_tx_data\[4\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.i_regbuf\[19\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[19\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[23\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_405 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_cycles.i_regbuf\[31\] i_tinyqv.cpu.i_core.i_cycles.reg_buf\[31\]
+ i_tinyqv.cpu.i_core.i_cycles.register\[3\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5170_ VGND VPWR _1925_ _1926_ _1924_ VPWR VGND sky130_fd_sc_hd__xnor2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.i_regbuf\[22\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[22\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[26\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4121_ VPWR VGND VGND VPWR i_tinyqv.cpu.data_addr\[2\] _0968_ _0967_ sky130_fd_sc_hd__nand2_1
X_4052_ VGND VPWR _0899_ _0784_ i_tinyqv.cpu.instr_data_start\[19\] _0898_ VPWR VGND
+ sky130_fd_sc_hd__and3_1
Xinput4 VGND VPWR net4 ui_in[2] VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7811_ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[30\] clknet_leaf_56_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[30\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4954_ VPWR VGND VPWR VGND _1727_ net97 _1732_ _0001_ sky130_fd_sc_hd__a21o_1
X_7742_ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[25\] clknet_leaf_55_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[25\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_3905_ VPWR VGND VPWR VGND i_tinyqv.cpu.i_core.i_registers.reg_access\[8\]\[1\] net27
+ _0757_ _0648_ i_tinyqv.cpu.i_core.i_registers.reg_access\[1\]\[1\] _0756_ sky130_fd_sc_hd__a221o_1
X_7673_ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[20\] clknet_leaf_59_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[20\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4885_ VGND VPWR VPWR VGND _1686_ _1184_ _1685_ i_tinyqv.cpu.i_core.i_registers.reg_access\[6\]\[0\]
+ sky130_fd_sc_hd__mux2_1
X_6624_ VGND VPWR i_tinyqv.cpu.was_early_branch _3017_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_3836_ _0688_ i_tinyqv.cpu.counter\[4\] VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_6555_ VPWR VGND VGND VPWR _2318_ _2952_ _2963_ _2964_ sky130_fd_sc_hd__o21a_1
XFILLER_0_14_121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_6_387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_6_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_3767_ VGND VPWR VGND VPWR _0619_ _0608_ _0614_ sky130_fd_sc_hd__nor2b_4
X_5506_ VPWR VGND _2216_ _2209_ i_uart_tx.cycle_counter\[6\] i_uart_tx.cycle_counter\[7\]
+ i_uart_tx.cycle_counter\[8\] VGND VPWR sky130_fd_sc_hd__a31o_1
X_6486_ VGND VPWR VPWR VGND _2903_ i_tinyqv.mem.q_ctrl.spi_in_buffer\[5\] _2897_ net133
+ sky130_fd_sc_hd__mux2_1
X_8225_ i_tinyqv.cpu.i_core.multiplier.accum\[8\] clknet_leaf_44_clk _0026_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5437_ VPWR VGND VPWR VGND _1679_ i_tinyqv.cpu.i_core.i_registers.rd\[3\] _2163_
+ _2164_ sky130_fd_sc_hd__a21oi_1
X_8156_ i_tinyqv.cpu.instr_data\[2\]\[5\] clknet_leaf_3_clk _0268_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5368_ VPWR VGND VPWR VGND _2087_ net211 _0840_ _0100_ _2101_ sky130_fd_sc_hd__a22o_1
X_8087_ gpio_out_sel\[6\] clknet_leaf_18_clk _0014_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4319_ VGND VPWR VGND VPWR net64 _0842_ _1166_ net45 sky130_fd_sc_hd__a21oi_4
X_5299_ _2048_ _0861_ _1752_ _1387_ _1031_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
X_7107_ VPWR VGND VPWR VGND _3308_ _2126_ _2143_ _3415_ sky130_fd_sc_hd__a21oi_1
X_7038_ VGND VPWR VPWR VGND _3350_ _3351_ _3349_ _3352_ sky130_fd_sc_hd__or3_2
Xi_tinyqv.cpu.i_core.i_cycles.i_regbuf\[5\] i_tinyqv.cpu.i_core.i_cycles.reg_buf\[5\]
+ i_tinyqv.cpu.i_core.cycle_count_wide\[5\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_157 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4670_ VGND VPWR VGND VPWR _1506_ i_tinyqv.cpu.instr_data\[0\]\[12\] _1504_ _1409_
+ _1505_ sky130_fd_sc_hd__o211a_1
X_6340_ VGND VPWR _0391_ _2781_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_614 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_6271_ VGND VPWR VPWR VGND _2745_ i_tinyqv.cpu.instr_data_in\[0\] _2744_ _2316_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_135 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.i_regbuf\[23\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[23\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[27\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_8010_ i_uart_rx.recieved_data\[3\] clknet_leaf_19_clk _0145_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.i_regbuf\[9\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[9\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[13\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5222_ VGND VPWR _1975_ _1976_ _1974_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_5153_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.multiplier.accum\[10\] _1910_ _1909_
+ sky130_fd_sc_hd__nand2_1
X_4104_ VGND VPWR VGND VPWR _0951_ _0927_ _0941_ i_tinyqv.cpu.i_core.cycle_count\[3\]
+ _0950_ sky130_fd_sc_hd__a211o_1
X_5084_ VGND VPWR VPWR VGND _1841_ _1844_ _1843_ sky130_fd_sc_hd__xor2_1
X_4035_ VPWR VGND _0882_ i_tinyqv.cpu.instr_data_start\[9\] VPWR VGND sky130_fd_sc_hd__buf_2
X_5986_ VGND VPWR _0262_ _2556_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4937_ VPWR VGND _1720_ i_tinyqv.cpu.instr_data_in\[14\] VPWR VGND sky130_fd_sc_hd__buf_2
X_7725_ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[8\] clknet_leaf_0_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[8\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XANTENNA_20 i_tinyqv.mem.q_ctrl.addr\[21\] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_0_62_514 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XANTENNA_31 i_tinyqv.cpu.i_core.imm_lo\[4\] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_7656_ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[3\] clknet_leaf_47_clk _0041_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4868_ VGND VPWR VPWR VGND _1676_ i_tinyqv.cpu.debug_rd\[1\] _1674_ i_tinyqv.cpu.i_core.i_registers.reg_access\[8\]\[1\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_205 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XANTENNA_42 i_tinyqv.cpu.i_core.imm_lo\[9\] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_6607_ VPWR VGND VGND VPWR _3002_ _3003_ _2061_ _0436_ sky130_fd_sc_hd__o21a_1
X_3819_ VGND VPWR VGND VPWR _0662_ _0663_ _0660_ _0671_ _0661_ sky130_fd_sc_hd__nor4b_2
X_4799_ VGND VPWR VGND VPWR _1634_ _1631_ _1633_ _0973_ _0752_ sky130_fd_sc_hd__a211o_1
X_7587_ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[30\] clknet_leaf_55_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[30\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6538_ VGND VPWR VPWR VGND _2949_ _2948_ _2920_ net13 sky130_fd_sc_hd__mux2_1
X_6469_ VPWR VGND VPWR VGND _2629_ i_tinyqv.cpu.i_core.i_shift.a\[28\] _2596_ _0409_
+ _2892_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_499 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_8208_ i_tinyqv.cpu.i_core.i_shift.a\[27\] clknet_leaf_40_clk _0320_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_8139_ i_tinyqv.cpu.data_addr\[14\] clknet_leaf_34_clk _0251_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.i_regbuf\[11\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[11\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[15\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.i_regbuf\[8\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[8\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[12\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_566 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_260 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xi_tinyqv.cpu.i_core.i_instrret.i_regbuf\[10\] i_tinyqv.cpu.i_core.i_instrret.reg_buf\[10\]
+ i_tinyqv.cpu.i_core.i_instrret.register\[14\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5840_ VGND VPWR VPWR VGND i_tinyqv.cpu.instr_write_offset\[2\] _1406_ _2460_ _2461_
+ sky130_fd_sc_hd__or3b_1
X_5771_ VGND VPWR _0194_ _2410_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_8490_ i_tinyqv.mem.q_ctrl.addr\[16\] clknet_leaf_32_clk _0588_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_4722_ VGND VPWR VGND VPWR i_tinyqv.cpu.data_read_n\[0\] i_tinyqv.cpu.data_read_n\[1\]
+ _1558_ net28 sky130_fd_sc_hd__a21oi_2
X_7510_ VGND VPWR _0599_ _3743_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7441_ VPWR VGND VPWR VGND _3681_ _0881_ _3010_ _3687_ sky130_fd_sc_hd__a21oi_1
X_4653_ VPWR VGND VGND VPWR _1489_ _1483_ _1488_ sky130_fd_sc_hd__or2_1
X_7372_ VGND VPWR _2682_ _3005_ _3629_ i_tinyqv.cpu.data_addr\[4\] VPWR VGND sky130_fd_sc_hd__o21ai_1
X_4584_ VGND VPWR VGND VPWR _1413_ _1419_ _1420_ _1409_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_4_655 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_6323_ VGND VPWR VPWR VGND _2773_ _2316_ _2772_ net279 sky130_fd_sc_hd__mux2_1
X_6254_ _2731_ _2708_ _2713_ _2722_ _2723_ _2728_ VPWR VGND VGND VPWR sky130_fd_sc_hd__o311a_1
X_5205_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.multiplier.accum\[12\] _1960_ _1959_
+ sky130_fd_sc_hd__nand2_1
X_6185_ VGND VPWR _0344_ _2673_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5136_ VGND VPWR VPWR VGND _1892_ _1894_ _1893_ sky130_fd_sc_hd__xor2_1
X_5067_ _1828_ _1803_ _1826_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
XFILLER_0_74_93 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4018_ VGND VPWR i_tinyqv.mem.qspi_data_byte_idx\[0\] _0868_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_5969_ VGND VPWR VPWR VGND _2545_ _2544_ _2501_ i_tinyqv.cpu.data_addr\[20\] sky130_fd_sc_hd__mux2_1
X_7708_ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[23\] clknet_leaf_59_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[23\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_385 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7639_ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[18\] clknet_leaf_46_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[18\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.i_regbuf\[23\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[23\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[27\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.i_regbuf\[12\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[12\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[16\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_419 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold109 net138 i_tinyqv.cpu.i_core.load_done VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7990_ i_uart_tx.cycle_counter\[9\] clknet_leaf_30_clk _0125_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_6941_ VGND VPWR VPWR VGND _0497_ _3274_ _3261_ _0691_ _3276_ net107 sky130_fd_sc_hd__a32o_1
X_6872_ VPWR VGND VPWR VGND _3240_ i_tinyqv.cpu.instr_fetch_stopped sky130_fd_sc_hd__inv_2
XFILLER_0_44_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_22_Left_103 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5823_ VPWR VGND VPWR VGND _2449_ _2448_ _2083_ _0207_ sky130_fd_sc_hd__a21oi_1
X_8542_ i_tinyqv.cpu.i_core.i_cycles.register\[15\] clknet_leaf_50_clk i_tinyqv.cpu.i_core.i_cycles.reg_buf\[15\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5754_ VPWR VGND VGND VPWR _2396_ _2198_ _2395_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_536 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5685_ VGND VPWR VGND VPWR _0174_ net97 _2330_ _2344_ _2299_ sky130_fd_sc_hd__o211a_1
X_4705_ VPWR VGND VPWR VGND _1541_ i_tinyqv.mem.qspi_write_done _1540_ sky130_fd_sc_hd__or2_2
X_8473_ i_tinyqv.cpu.additional_mem_ops\[2\] clknet_leaf_6_clk _0571_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_7424_ VGND VPWR VGND VPWR _3673_ _3632_ _3671_ _3672_ _2681_ sky130_fd_sc_hd__o211a_1
X_4636_ VGND VPWR VGND VPWR _1472_ i_tinyqv.cpu.instr_data\[0\]\[13\] _1414_ _1408_
+ _1471_ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_539 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_4_485 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7355_ VGND VPWR VPWR VGND _0571_ _3615_ _2049_ net154 _3616_ _3359_ sky130_fd_sc_hd__a32o_1
X_6306_ VGND VPWR _0375_ _2763_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_31_Left_112 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4567_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.mie\[19\] _1403_ _0991_ sky130_fd_sc_hd__nand2_1
X_7286_ VGND VPWR _0557_ _3561_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4498_ VPWR VGND VGND VPWR i_tinyqv.cpu.instr_data_start\[14\] _0895_ _1337_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_296 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_40_583 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6237_ VPWR VGND VGND VPWR _1060_ _2716_ _1880_ sky130_fd_sc_hd__nand2_1
X_6168_ VGND VPWR _0336_ _2664_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5119_ VPWR VGND VGND VPWR _1859_ _1877_ _1860_ sky130_fd_sc_hd__nand2_1
X_6099_ VGND VPWR _0314_ _2617_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_40_Left_121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5470_ VGND VPWR VPWR VGND _2191_ i_uart_tx.data_to_send\[6\] _2177_ i_uart_tx.data_to_send\[5\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_4421_ VPWR VGND VGND VPWR _1149_ _1087_ _1264_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_4352_ VPWR VGND VPWR VGND _0944_ i_tinyqv.cpu.i_core.mip\[17\] _0943_ _1195_ i_tinyqv.cpu.i_core.mie\[17\]
+ sky130_fd_sc_hd__a22o_1
X_7140_ VGND VPWR VGND VPWR _3445_ _3300_ _3444_ _3298_ _2120_ sky130_fd_sc_hd__o211a_1
X_4283_ VGND VPWR VPWR VGND _1130_ _1093_ _1103_ _1072_ sky130_fd_sc_hd__mux2_1
X_7071_ VPWR VGND VPWR VGND i_tinyqv.cpu.instr_data\[3\]\[5\] _3369_ _3383_ _3370_
+ i_tinyqv.cpu.instr_data\[2\]\[5\] _3372_ sky130_fd_sc_hd__a221o_1
X_6022_ VGND VPWR VPWR VGND _2577_ i_tinyqv.cpu.instr_data\[2\]\[15\] _2562_ _1721_
+ sky130_fd_sc_hd__mux2_1
X_7973_ i_uart_tx.data_to_send\[0\] clknet_leaf_29_clk _0108_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_6924_ VGND VPWR VPWR VGND _0485_ _3265_ _3261_ _1589_ _3271_ net149 sky130_fd_sc_hd__a32o_1
X_6855_ VPWR VGND VGND VPWR i_tinyqv.cpu.instr_data_start\[22\] i_tinyqv.cpu.imm\[22\]
+ _3225_ sky130_fd_sc_hd__nor2_1
X_6786_ VGND VPWR VGND VPWR _3163_ _3159_ _3162_ _3051_ _3029_ sky130_fd_sc_hd__a211o_1
XFILLER_0_9_566 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_3998_ VGND VPWR _0653_ i_tinyqv.cpu.is_alu_reg _0849_ i_tinyqv.cpu.is_alu_imm VPWR
+ VGND sky130_fd_sc_hd__o21ai_2
X_5806_ VPWR VGND VPWR VGND _0907_ _0752_ _2435_ _2434_ _2433_ sky130_fd_sc_hd__or4bb_1
X_5737_ VPWR VGND VGND VPWR _2381_ i_spi.clock_divider\[1\] i_spi.clock_count\[1\]
+ sky130_fd_sc_hd__or2_1
X_8525_ i_tinyqv.cpu.i_core.i_instrret.register\[31\] clknet_leaf_47_clk i_tinyqv.cpu.i_core.i_instrret.reg_buf\[31\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_8456_ i_tinyqv.cpu.alu_op\[2\] clknet_leaf_39_clk _0554_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5668_ VPWR VGND VPWR VGND _0989_ _2328_ _0995_ _2329_ sky130_fd_sc_hd__or3_1
X_7407_ VGND VPWR VGND VPWR _3659_ i_tinyqv.cpu.data_addr\[9\] _3012_ _3004_ _3658_
+ sky130_fd_sc_hd__o211a_1
X_5599_ VPWR VGND VPWR VGND _2281_ _2238_ _2280_ sky130_fd_sc_hd__or2_2
X_8387_ i_tinyqv.cpu.data_out\[12\] clknet_leaf_19_clk _0485_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.i_regbuf\[26\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[26\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[30\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4619_ VGND VPWR VPWR VGND _1409_ _1454_ _1453_ _1455_ sky130_fd_sc_hd__mux2_2
X_7338_ VGND VPWR VPWR VGND _3605_ _0661_ _2153_ _3604_ sky130_fd_sc_hd__mux2_1
X_7269_ VGND VPWR _0554_ _3547_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_406 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_55_439 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_3_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_35_163 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_51_634 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_50_111 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4970_ VPWR VGND VGND VPWR _1742_ net14 _1725_ sky130_fd_sc_hd__nand2_2
X_3921_ VGND VPWR VGND VPWR i_tinyqv.cpu.imm\[21\] i_tinyqv.cpu.imm\[17\] _0608_ i_tinyqv.cpu.imm\[29\]
+ i_tinyqv.cpu.imm\[25\] _0614_ _0773_ sky130_fd_sc_hd__mux4_1
X_6640_ VGND VPWR VGND VPWR _3031_ _2995_ _3002_ _1339_ _3029_ sky130_fd_sc_hd__a211o_1
X_3852_ VPWR VGND VPWR VGND i_tinyqv.cpu.i_core.imm_lo\[0\] _0615_ _0704_ _0620_ i_tinyqv.cpu.i_core.imm_lo\[8\]
+ i_tinyqv.cpu.counter\[4\] sky130_fd_sc_hd__a221o_1
X_6571_ VGND VPWR _0426_ _2977_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5522_ VGND VPWR _2228_ _2226_ _2181_ _2227_ VPWR VGND sky130_fd_sc_hd__and3_1
X_3783_ VPWR VGND VPWR VGND net321 i_tinyqv.cpu.i_core.i_registers.reg_access\[15\]\[3\]
+ _0633_ _0635_ i_tinyqv.cpu.i_core.i_registers.reg_access\[8\]\[3\] sky130_fd_sc_hd__a22o_1
X_8310_ i_tinyqv.cpu.i_core.i_shift.a\[28\] clknet_leaf_39_clk _0409_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
X_5453_ _0991_ _2179_ _0997_ _1557_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_8241_ i_tinyqv.cpu.i_core.mepc\[12\] clknet_leaf_35_clk _0341_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_4404_ VPWR VGND VGND VPWR _1247_ _1169_ _1246_ sky130_fd_sc_hd__or2_1
X_5384_ VPWR VGND _0102_ _2115_ _2114_ _2057_ _2083_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_8172_ i_tinyqv.cpu.instr_data\[1\]\[7\] clknet_leaf_10_clk _0284_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_4335_ VGND VPWR VPWR VGND _1182_ _1169_ _1168_ _0846_ _1170_ _1181_ sky130_fd_sc_hd__a32o_1
X_7123_ VPWR VGND VGND VPWR _1478_ _3352_ _1510_ _3430_ sky130_fd_sc_hd__o21a_1
X_4266_ VGND VPWR VPWR VGND _1113_ i_tinyqv.cpu.i_core.i_shift.a\[14\] _1028_ i_tinyqv.cpu.i_core.i_shift.a\[17\]
+ sky130_fd_sc_hd__mux2_1
X_7054_ VPWR VGND VGND VPWR _1422_ _3367_ _1432_ sky130_fd_sc_hd__nand2_1
X_4197_ VPWR VGND VPWR VGND _1039_ i_tinyqv.cpu.i_core.i_shift.b\[3\] _1043_ _1044_
+ sky130_fd_sc_hd__a21o_1
X_6005_ VGND VPWR _0269_ _2568_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7956_ i_tinyqv.cpu.i_core.time_hi\[2\] clknet_leaf_51_clk _0094_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_6907_ VPWR VGND _3263_ _3262_ _1026_ VPWR VGND sky130_fd_sc_hd__and2_1
X_7887_ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[10\] clknet_leaf_5_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[10\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6838_ VGND VPWR VGND VPWR _3208_ _3210_ _3209_ sky130_fd_sc_hd__or2b_1
X_6769_ VPWR VGND VGND VPWR i_tinyqv.cpu.instr_data_start\[14\] i_tinyqv.cpu.imm\[14\]
+ _3147_ sky130_fd_sc_hd__nor2_1
X_8508_ i_tinyqv.cpu.i_core.i_instrret.register\[14\] clknet_leaf_49_clk i_tinyqv.cpu.i_core.i_instrret.reg_buf\[14\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_612 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.i_regbuf\[27\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[27\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[31\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_8439_ i_tinyqv.cpu.imm\[17\] clknet_leaf_22_clk _0537_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_13_380 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold270 net299 i_tinyqv.cpu.data_addr\[5\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 net310 i_tinyqv.mem.q_ctrl.addr\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.i_regbuf\[30\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[30\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[2\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.i_regbuf\[26\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[26\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[30\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_539 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xi_tinyqv.cpu.i_core.i_cycles.i_regbuf\[24\] i_tinyqv.cpu.i_core.i_cycles.reg_buf\[24\]
+ i_tinyqv.cpu.i_core.i_cycles.register\[28\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4120_ VPWR VGND VGND VPWR _0966_ _0961_ i_tinyqv.cpu.data_addr\[5\] _0967_ sky130_fd_sc_hd__nor3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.i_regbuf\[15\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[15\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[19\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4051_ VPWR VGND _0898_ _0897_ i_tinyqv.cpu.instr_data_start\[17\] VPWR VGND sky130_fd_sc_hd__and2_1
Xinput5 VPWR VGND net5 ui_in[3] VPWR VGND sky130_fd_sc_hd__buf_2
X_7810_ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[29\] clknet_leaf_57_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[29\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4953_ VGND VPWR _1732_ gpio_out\[1\] _1729_ _1730_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_59_575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_7741_ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[24\] clknet_leaf_59_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[24\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_74 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_7672_ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[19\] clknet_leaf_46_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[19\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_3904_ VPWR VGND VPWR VGND i_tinyqv.cpu.i_core.i_registers.reg_access\[2\]\[1\] net26
+ _0756_ _0646_ i_tinyqv.cpu.i_core.i_registers.reg_access\[10\]\[1\] _0755_ sky130_fd_sc_hd__a221o_1
X_6623_ VPWR VGND VGND VPWR _3016_ _0884_ i_tinyqv.cpu.instr_write_offset\[3\] sky130_fd_sc_hd__or2_1
X_4884_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_registers.rd\[3\] _1188_ _1641_
+ i_tinyqv.cpu.i_core.i_registers.rd\[2\] _1685_ sky130_fd_sc_hd__and4b_2
XFILLER_0_46_258 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_3835_ VPWR VGND VGND VPWR _0686_ _0687_ _0673_ sky130_fd_sc_hd__nor2_2
X_6554_ VGND VPWR VGND VPWR _2963_ _2960_ _2962_ _2914_ _2956_ sky130_fd_sc_hd__a211o_1
X_3766_ VPWR VGND VPWR VGND _0617_ i_tinyqv.cpu.instr_data_start\[3\] _0615_ _0618_
+ i_tinyqv.cpu.instr_data_start\[15\] sky130_fd_sc_hd__a22o_1
X_6485_ VGND VPWR _0415_ net168 VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5505_ VGND VPWR _2215_ net157 net170 _2212_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_72_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_8224_ i_tinyqv.cpu.i_core.multiplier.accum\[7\] clknet_leaf_44_clk _0025_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5436_ VGND VPWR _1679_ _2149_ _2163_ i_tinyqv.cpu.i_core.i_registers.rd\[3\] VPWR
+ VGND sky130_fd_sc_hd__o21ai_1
X_5367_ VPWR VGND VPWR VGND _2099_ _0623_ _2056_ _2101_ _2100_ sky130_fd_sc_hd__a22o_1
X_8155_ i_tinyqv.cpu.instr_data\[2\]\[4\] clknet_leaf_10_clk _0267_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_8086_ gpio_out_sel\[5\] clknet_leaf_18_clk _0013_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4318_ VGND VPWR _1165_ _1125_ _1123_ _1164_ VPWR VGND sky130_fd_sc_hd__and3_1
X_5298_ VPWR VGND VPWR VGND _1026_ net138 _2047_ _0084_ sky130_fd_sc_hd__a21o_1
X_7106_ VGND VPWR _0524_ _3414_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4249_ VGND VPWR VPWR VGND _1096_ i_tinyqv.cpu.i_core.i_shift.a\[26\] _1036_ i_tinyqv.cpu.i_core.i_shift.a\[5\]
+ sky130_fd_sc_hd__mux2_1
X_7037_ _2123_ _3351_ _1426_ _3322_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_7939_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[30\] clknet_leaf_49_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[30\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_203 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_37_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_65_545 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_18_472 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_21_659 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.i_regbuf\[31\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[31\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[3\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_78_Left_159 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_51_250 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6270_ VGND VPWR _2743_ _2744_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_5221_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[11\] _1975_ _1880_ sky130_fd_sc_hd__nand2_1
X_5152_ VPWR VGND _1909_ _1908_ _1907_ VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_20_692 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.i_regbuf\[16\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[16\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[20\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4103_ VPWR VGND VPWR VGND i_tinyqv.cpu.i_core.mip\[16\] _0943_ _0950_ _0944_ i_tinyqv.cpu.i_core.mie\[16\]
+ _0949_ sky130_fd_sc_hd__a221o_1
X_5083_ VPWR VGND VPWR VGND _1816_ i_tinyqv.cpu.i_core.multiplier.accum\[6\] _1842_
+ _1843_ sky130_fd_sc_hd__a21o_1
XFILLER_0_47_74 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4034_ VPWR VGND _0881_ i_tinyqv.cpu.instr_data_start\[15\] VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_0_63_40 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_66_309 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7724_ i_tinyqv.cpu.i_core.i_registers.reg_access\[9\]\[3\] clknet_leaf_53_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[7\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5985_ VPWR VGND _2556_ _2555_ _2079_ VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_74_342 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4936_ VGND VPWR VGND VPWR _1711_ _1717_ _1719_ uio_out[2] _1718_ sky130_fd_sc_hd__a211o_4
XANTENNA_21 i_tinyqv.mem.q_ctrl.addr\[21\] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_10 _3068_ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_7655_ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[2\] clknet_leaf_47_clk _0040_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4867_ VGND VPWR _0074_ _1675_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XANTENNA_32 i_tinyqv.cpu.i_core.is_interrupt VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_43 i_tinyqv.cpu.i_core.imm_lo\[9\] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_6606_ _3003_ _1524_ _2995_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
XFILLER_0_6_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7586_ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[29\] clknet_leaf_58_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[29\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_3818_ VPWR VGND VGND VPWR _0661_ _0670_ _0660_ sky130_fd_sc_hd__nor2_2
XFILLER_0_34_217 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6537_ VGND VPWR VPWR VGND _2948_ i_tinyqv.mem.q_ctrl.spi_in_buffer\[3\] _2918_ i_tinyqv.mem.q_ctrl.spi_in_buffer\[7\]
+ sky130_fd_sc_hd__mux2_1
X_4798_ VGND VPWR VGND VPWR _1633_ _0970_ _0969_ _1632_ _0968_ sky130_fd_sc_hd__o211a_1
X_6468_ VGND VPWR _1124_ _2891_ _2892_ _1312_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_6399_ VPWR VGND VGND VPWR _1540_ _2836_ _2787_ sky130_fd_sc_hd__nand2_1
X_8207_ i_tinyqv.cpu.i_core.i_shift.a\[26\] clknet_leaf_40_clk _0319_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5419_ _0863_ _2149_ _0837_ _1440_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_8138_ i_tinyqv.cpu.data_addr\[13\] clknet_leaf_34_clk _0250_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_8069_ i_spi.clock_divider\[1\] clknet_leaf_27_clk _0204_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xmax_cap23 VGND VPWR net23 _0714_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_401 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_68_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_5770_ VPWR VGND _2410_ _2409_ _2221_ VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_29_545 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_4721_ VGND VPWR VGND VPWR i_tinyqv.cpu.data_write_n\[0\] net28 _1557_ i_tinyqv.cpu.data_write_n\[1\]
+ sky130_fd_sc_hd__a21oi_4
XFILLER_0_29_567 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_56_397 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7440_ VPWR VGND VGND VPWR _3686_ _0881_ _3681_ sky130_fd_sc_hd__or2_1
X_4652_ VPWR VGND VGND VPWR _1488_ _1426_ _1487_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_634 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_7371_ VPWR VGND VGND VPWR _3626_ _3627_ _3045_ _3239_ _3628_ _2681_ sky130_fd_sc_hd__o221a_1
X_4583_ VGND VPWR VGND VPWR _1419_ i_tinyqv.cpu.instr_data\[1\]\[0\] _1414_ _1416_
+ _1418_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_645 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_40_710 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6322_ VGND VPWR _2771_ _2772_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_294 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_6253_ VPWR VGND VGND VPWR _2696_ _2730_ _2726_ sky130_fd_sc_hd__nand2_1
X_5204_ VPWR VGND _1959_ _1958_ _1957_ VPWR VGND sky130_fd_sc_hd__and2_1
X_6184_ VGND VPWR VPWR VGND _2673_ i_tinyqv.cpu.i_core.mepc\[19\] _2667_ i_tinyqv.cpu.i_core.mepc\[15\]
+ sky130_fd_sc_hd__mux2_1
X_5135_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[8\] _1893_ _1845_ sky130_fd_sc_hd__nand2_1
X_5066_ _1803_ _1825_ _1827_ _1826_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_4017_ VGND VPWR _0866_ _0867_ _0864_ VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_640 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.i_regbuf\[20\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[20\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[24\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5968_ VGND VPWR VPWR VGND _2544_ i_tinyqv.cpu.i_core.mepc\[20\] _2106_ i_tinyqv.cpu.i_core.i_shift.a\[24\]
+ sky130_fd_sc_hd__mux2_1
X_7707_ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[22\] clknet_leaf_52_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[22\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4919_ VGND VPWR VPWR VGND _1705_ _1638_ _1701_ i_tinyqv.cpu.i_core.i_registers.reg_access\[1\]\[3\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_353 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5899_ VGND VPWR VPWR VGND _2497_ _2496_ _2399_ i_spi.data\[6\] sky130_fd_sc_hd__mux2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.i_regbuf\[6\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[6\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[10\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7638_ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[17\] clknet_leaf_55_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[17\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7569_ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[12\] clknet_leaf_58_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[12\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.i_regbuf\[16\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[16\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[20\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.i_regbuf\[4\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[4\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[8\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_39 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_22_710 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_6940_ VPWR VGND VGND VPWR _3276_ _0630_ _0854_ sky130_fd_sc_hd__or2_1
X_6871_ VGND VPWR _1437_ _3239_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_640 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5822_ VPWR VGND VGND VPWR _0944_ _2449_ _2103_ sky130_fd_sc_hd__nand2_1
X_5753_ VPWR VGND VGND VPWR _2392_ _2394_ _2395_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_8541_ i_tinyqv.cpu.i_core.i_cycles.register\[14\] clknet_leaf_5_clk i_tinyqv.cpu.i_core.i_cycles.reg_buf\[14\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4704_ VGND VPWR _1539_ _1540_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_5684_ VGND VPWR VGND VPWR _2344_ _2336_ _2341_ net233 _2343_ sky130_fd_sc_hd__a211o_1
X_8472_ i_tinyqv.cpu.additional_mem_ops\[1\] clknet_leaf_6_clk _0570_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_7423_ VPWR VGND VGND VPWR _3632_ _3672_ _3129_ sky130_fd_sc_hd__nand2_1
X_4635_ VPWR VGND VGND VPWR _1471_ i_tinyqv.cpu.instr_data\[2\]\[13\] _1417_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_710 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_8_75 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_7354_ VPWR VGND VPWR VGND _3351_ _1501_ _2143_ _3616_ _1491_ sky130_fd_sc_hd__a22o_1
X_4566_ VPWR VGND VPWR VGND _1228_ i_tinyqv.cpu.i_core.mie\[18\] _1401_ _1402_ sky130_fd_sc_hd__a21oi_1
X_6305_ VGND VPWR VPWR VGND _2763_ _2316_ _2762_ net280 sky130_fd_sc_hd__mux2_1
XFILLER_0_12_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7285_ VGND VPWR VPWR VGND _3561_ _3560_ _3395_ i_tinyqv.cpu.i_core.mem_op\[1\] sky130_fd_sc_hd__mux2_1
X_4497_ VPWR VGND VGND VPWR _0610_ _1336_ _1335_ sky130_fd_sc_hd__nand2_1
X_6236_ VPWR VGND VGND VPWR _2715_ _2700_ _2701_ sky130_fd_sc_hd__or2_1
X_6167_ VGND VPWR VPWR VGND _2664_ i_tinyqv.cpu.i_core.mepc\[11\] _2656_ i_tinyqv.cpu.i_core.mepc\[7\]
+ sky130_fd_sc_hd__mux2_1
X_5118_ VGND VPWR _0022_ _1876_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6098_ VGND VPWR VPWR VGND _2617_ i_tinyqv.cpu.i_core.i_shift.a\[21\] _2595_ i_tinyqv.cpu.i_core.i_shift.a\[25\]
+ sky130_fd_sc_hd__mux2_1
X_5049_ VPWR VGND VGND VPWR _1808_ _1810_ _1809_ sky130_fd_sc_hd__nand2_1
Xclone11 VGND VPWR _1398_ net40 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.i_regbuf\[20\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[20\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[24\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_23 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_45_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_26_312 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_54_665 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4420_ VPWR VGND VGND VPWR _1092_ _1263_ _1262_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_337 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4351_ VGND VPWR _1194_ uo_out[5] VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_4282_ VPWR VGND VGND VPWR _1092_ _1129_ _1128_ sky130_fd_sc_hd__nand2_1
X_7070_ VGND VPWR VPWR VGND _3377_ _3355_ _3381_ _3382_ sky130_fd_sc_hd__or3b_1
X_6021_ VGND VPWR _0277_ _2576_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7972_ i_tinyqv.cpu.i_core.i_cycles.rstn clknet_leaf_17_clk i_debug_uart_tx.resetn
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_55_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6923_ VGND VPWR VPWR VGND _0724_ _0854_ _0956_ _3271_ sky130_fd_sc_hd__or3_2
X_6854_ VPWR VGND VPWR VGND _3215_ _3224_ _3216_ _3218_ sky130_fd_sc_hd__a21boi_1
X_6785_ VPWR VGND VGND VPWR _2993_ _3161_ _3162_ sky130_fd_sc_hd__nor2_1
X_3997_ VPWR VGND VGND VPWR _0842_ _0847_ _0848_ sky130_fd_sc_hd__nor2_1
X_5805_ VPWR VGND VGND VPWR _2434_ _0920_ _0944_ sky130_fd_sc_hd__nand2_2
X_5736_ VPWR VGND VGND VPWR i_spi.clock_divider\[1\] _2380_ i_spi.clock_count\[1\]
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_492 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_9_589 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_8524_ i_tinyqv.cpu.i_core.i_instrret.register\[30\] clknet_leaf_50_clk i_tinyqv.cpu.i_core.i_instrret.reg_buf\[30\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5667_ VPWR VGND VGND VPWR _0984_ _0987_ _2328_ _1557_ sky130_fd_sc_hd__nand3_1
X_8455_ i_tinyqv.cpu.alu_op\[1\] clknet_leaf_38_clk _0553_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7406_ VPWR VGND VPWR VGND _3632_ _3099_ _3658_ _3656_ _3657_ _2877_ sky130_fd_sc_hd__a221o_1
X_4618_ VGND VPWR VPWR VGND _1454_ i_tinyqv.cpu.instr_data\[2\]\[6\] _1414_ i_tinyqv.cpu.instr_data\[0\]\[6\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5598_ VGND VPWR _1227_ i_uart_rx.fsm_state\[0\] _2280_ _2239_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_8386_ i_tinyqv.cpu.data_out\[11\] clknet_leaf_26_clk _0484_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_4549_ VPWR VGND VPWR VGND _1385_ i_tinyqv.cpu.data_continue sky130_fd_sc_hd__inv_2
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.i_regbuf\[19\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[19\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[23\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7337_ VGND VPWR VPWR VGND _3604_ _3603_ _2147_ _3601_ sky130_fd_sc_hd__mux2_1
X_7268_ VGND VPWR VPWR VGND _3547_ _3546_ _3395_ _1030_ sky130_fd_sc_hd__mux2_1
X_6219_ VPWR VGND VGND VPWR _2695_ _2026_ _2699_ _2697_ sky130_fd_sc_hd__nand3_1
X_7199_ VGND VPWR VGND VPWR _3495_ i_tinyqv.cpu.instr_data\[2\]\[1\] _1432_ _1423_
+ _3489_ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_51_613 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_63_484 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_35_175 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_50_156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_3920_ VPWR VGND VGND VPWR _0768_ _0766_ _0772_ _0771_ sky130_fd_sc_hd__nor3_4
X_3851_ VPWR VGND VPWR VGND _0619_ i_tinyqv.cpu.imm\[12\] _0617_ _0703_ i_tinyqv.cpu.i_core.imm_lo\[4\]
+ sky130_fd_sc_hd__a22o_1
X_6570_ VGND VPWR VPWR VGND _2977_ _1721_ _2925_ _2976_ sky130_fd_sc_hd__mux2_1
X_3782_ VPWR VGND VGND VPWR _0626_ _0625_ _0634_ _0624_ _0627_ sky130_fd_sc_hd__nor4b_1
X_5521_ VPWR VGND VPWR VGND _2225_ i_uart_tx.fsm_state\[0\] i_uart_tx.fsm_state\[1\]
+ _2227_ sky130_fd_sc_hd__a21o_1
XFILLER_0_42_624 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_8240_ i_tinyqv.cpu.i_core.mepc\[11\] clknet_leaf_35_clk _0340_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_5452_ VGND VPWR VPWR VGND _2178_ i_uart_tx.data_to_send\[1\] _2177_ i_uart_tx.data_to_send\[0\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_359 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_42_679 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_220 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4403_ VPWR VGND VGND VPWR _1246_ _1244_ _1245_ sky130_fd_sc_hd__or2_1
X_8171_ i_tinyqv.cpu.instr_data\[1\]\[6\] clknet_leaf_10_clk _0283_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5383_ VPWR VGND VGND VPWR _2115_ net262 _1393_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_554 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4334_ VGND VPWR VGND VPWR _1181_ _1174_ _1176_ _1172_ _1180_ sky130_fd_sc_hd__a211o_1
X_7122_ VGND VPWR VGND VPWR _2133_ _3428_ _3329_ _3429_ _1460_ sky130_fd_sc_hd__a2bb2o_1
X_7053_ VGND VPWR _3365_ _3366_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_4265_ VGND VPWR VPWR VGND _1112_ _1111_ _1103_ _1110_ sky130_fd_sc_hd__mux2_1
X_6004_ VGND VPWR VPWR VGND _2568_ i_tinyqv.cpu.instr_data\[2\]\[6\] _2563_ i_tinyqv.cpu.instr_data_in\[6\]
+ sky130_fd_sc_hd__mux2_1
X_4196_ VPWR VGND VGND VPWR _1040_ _1042_ _1043_ sky130_fd_sc_hd__nor2_1
X_7955_ i_tinyqv.cpu.i_core.time_hi\[1\] clknet_leaf_51_clk _0093_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_6906_ VPWR VGND VGND VPWR _0956_ _3262_ _0612_ sky130_fd_sc_hd__nand2_1
X_7886_ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[9\] clknet_leaf_5_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[9\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6837_ VPWR VGND VGND VPWR i_tinyqv.cpu.instr_data_start\[20\] _3209_ i_tinyqv.cpu.imm\[20\]
+ sky130_fd_sc_hd__nand2_1
X_6768_ _3146_ _3138_ _3126_ _3139_ _3136_ VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_8507_ i_tinyqv.cpu.i_core.i_instrret.register\[13\] clknet_leaf_45_clk i_tinyqv.cpu.i_core.i_instrret.reg_buf\[13\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_462 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_5719_ VPWR VGND VGND VPWR i_debug_uart_tx.fsm_state\[3\] _2367_ i_debug_uart_tx.fsm_state\[1\]
+ sky130_fd_sc_hd__nand2_1
X_6699_ VPWR VGND VPWR VGND _3083_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[16\]
+ sky130_fd_sc_hd__inv_2
X_8438_ i_tinyqv.cpu.imm\[16\] clknet_leaf_8_clk _0536_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_8369_ i_tinyqv.cpu.data_write_n\[1\] clknet_leaf_21_clk _0468_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_32_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold260 net289 i_tinyqv.mem.q_ctrl.spi_flash_select VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 net300 i_tinyqv.cpu.data_addr\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 net311 i_tinyqv.mem.q_ctrl.spi_ram_b_select VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.i_regbuf\[23\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[23\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[27\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_11_68 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.i_regbuf\[19\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[19\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[23\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_cycles.i_regbuf\[17\] i_tinyqv.cpu.i_core.i_cycles.reg_buf\[17\]
+ i_tinyqv.cpu.i_core.i_cycles.register\[21\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4050_ VGND VPWR _0897_ _0881_ i_tinyqv.cpu.instr_data_start\[16\] _0896_ VPWR VGND
+ sky130_fd_sc_hd__and3_1
Xinput6 VGND VPWR ui_in[4] net6 VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_4952_ VPWR VGND VPWR VGND _1727_ net117 _1731_ _0000_ sky130_fd_sc_hd__a21o_1
X_7740_ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[23\] clknet_leaf_53_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[23\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7671_ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[18\] clknet_leaf_58_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[18\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_3903_ VPWR VGND VPWR VGND net46 i_tinyqv.cpu.i_core.i_registers.reg_access\[12\]\[1\]
+ net75 _0755_ i_tinyqv.cpu.i_core.i_registers.reg_access\[14\]\[1\] sky130_fd_sc_hd__a22o_1
X_4883_ VGND VPWR _0073_ _1684_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6622_ VPWR VGND VPWR VGND _3015_ net126 _3009_ _0439_ _3005_ sky130_fd_sc_hd__a22o_1
X_3834_ VGND VPWR VPWR VGND _0685_ _0682_ _0679_ _0676_ _0686_ sky130_fd_sc_hd__or4_4
X_6553_ VGND VPWR VGND VPWR _2962_ i_tinyqv.cpu.data_out\[13\] _2912_ _2929_ _2961_
+ sky130_fd_sc_hd__o211a_1
X_3765_ VPWR VGND _0617_ _0616_ VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_0_14_101 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_15_624 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_484 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_42_421 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5504_ VPWR VGND VPWR VGND _2212_ net157 _2214_ _0123_ sky130_fd_sc_hd__a21oi_1
X_6484_ VGND VPWR VPWR VGND _2902_ i_tinyqv.mem.q_ctrl.spi_in_buffer\[4\] _2897_ net167
+ sky130_fd_sc_hd__mux2_1
X_8223_ i_tinyqv.cpu.i_core.multiplier.accum\[6\] clknet_leaf_44_clk _0024_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5435_ VPWR VGND VPWR VGND _2153_ i_tinyqv.cpu.i_core.i_registers.rd\[2\] _2162_
+ _0106_ sky130_fd_sc_hd__a21o_1
X_8154_ i_tinyqv.cpu.instr_data\[2\]\[3\] clknet_leaf_11_clk _0266_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5366_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.mepc\[3\] net18 _1395_ _2100_ sky130_fd_sc_hd__o21a_1
X_8085_ gpio_out_sel\[4\] clknet_leaf_18_clk _0012_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_395 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_4317_ VPWR VGND VGND VPWR _0843_ _1164_ _1163_ sky130_fd_sc_hd__nand2_1
X_5297_ VGND VPWR _2047_ i_tinyqv.cpu.i_core.cycle\[1\] i_tinyqv.cpu.data_ready_core
+ _0744_ VPWR VGND sky130_fd_sc_hd__and3_1
X_7105_ VGND VPWR VPWR VGND _3414_ _3413_ _3396_ i_tinyqv.cpu.i_core.imm_lo\[4\] sky130_fd_sc_hd__mux2_1
X_4248_ VGND VPWR VPWR VGND _1095_ _1094_ _1083_ _1093_ sky130_fd_sc_hd__mux2_1
X_7036_ VPWR VGND _3350_ _3322_ _1468_ VPWR VGND sky130_fd_sc_hd__and2_1
X_4179_ VGND VPWR _0946_ _1026_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_7938_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[29\] clknet_leaf_50_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[29\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7869_ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[24\] clknet_leaf_48_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[24\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_3__f_clk VGND VPWR VGND VPWR clknet_0_clk clknet_3_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_14_Right_14 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_33_454 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_23_Right_23 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.i_regbuf\[24\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[24\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[28\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_32_Right_32 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_24_421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_24_432 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5220_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[10\] _1974_ _1813_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_41_Right_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5151_ VPWR VGND VGND VPWR _1908_ _1905_ _1906_ sky130_fd_sc_hd__or2_1
X_5082_ VPWR VGND _1842_ _1815_ _1812_ VPWR VGND sky130_fd_sc_hd__and2_1
X_4102_ VPWR VGND VPWR VGND _0948_ i_tinyqv.cpu.i_core.mcause\[0\] _0947_ _0949_ i_tinyqv.cpu.i_core.mepc\[0\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_42 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4033_ VGND VPWR _0879_ _0880_ VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_0_79_605 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_50_Right_50 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7723_ i_tinyqv.cpu.i_core.i_registers.reg_access\[9\]\[2\] clknet_leaf_1_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[6\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5984_ VPWR VGND VPWR VGND _2552_ i_tinyqv.cpu.data_addr\[25\] _1758_ _2555_ i_tinyqv.cpu.i_core.i_shift.a\[29\]
+ sky130_fd_sc_hd__a22o_1
X_4935_ VPWR VGND VGND VPWR _1706_ _1708_ _1714_ _1719_ sky130_fd_sc_hd__o21a_1
XANTENNA_11 i_tinyqv.cpu.data_addr\[24\] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_22 i_tinyqv.mem.q_ctrl.addr\[21\] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_0_7_621 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_7654_ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[1\] clknet_leaf_55_clk _0039_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4866_ VGND VPWR VPWR VGND _1675_ i_tinyqv.cpu.debug_rd\[0\] _1674_ i_tinyqv.cpu.i_core.i_registers.reg_access\[8\]\[0\]
+ sky130_fd_sc_hd__mux2_1
X_4797_ VPWR VGND VPWR VGND i_tinyqv.mem.data_from_read\[19\] _0689_ _1632_ _0748_
+ i_tinyqv.mem.data_from_read\[23\] _0865_ sky130_fd_sc_hd__a221o_1
X_6605_ VPWR VGND VPWR VGND _3001_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[10\]
+ _2987_ _3002_ _2993_ sky130_fd_sc_hd__a22o_1
XANTENNA_44 i_tinyqv.cpu.i_core.imm_lo\[9\] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.i_regbuf\[12\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[12\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[16\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7585_ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[28\] clknet_leaf_59_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[28\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_3817_ VGND VPWR VPWR VGND _0669_ _0667_ _0666_ i_tinyqv.cpu.i_core.i_registers.reg_access\[10\]\[3\]
+ _0668_ i_tinyqv.cpu.i_core.i_registers.reg_access\[14\]\[3\] sky130_fd_sc_hd__a32o_1
XANTENNA_33 i_tinyqv.cpu.i_core.mepc\[3\] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_6536_ VGND VPWR VPWR VGND _2947_ _2946_ _2916_ net13 sky130_fd_sc_hd__mux2_1
XFILLER_0_6_175 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_6467_ VGND VPWR VGND VPWR _2891_ _2625_ _2890_ _2640_ _0845_ sky130_fd_sc_hd__a211o_1
X_6398_ VGND VPWR _0395_ _2835_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_381 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5418_ VGND VPWR VPWR VGND _2148_ _2145_ _2147_ _1640_ sky130_fd_sc_hd__mux2_1
X_8206_ i_tinyqv.cpu.i_core.i_shift.a\[25\] clknet_leaf_40_clk _0318_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5349_ VGND VPWR _0096_ _2086_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8137_ i_tinyqv.cpu.data_addr\[12\] clknet_leaf_34_clk _0249_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_8068_ i_spi.clock_divider\[0\] clknet_leaf_27_clk net163 VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7019_ _3336_ _2119_ _1476_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
Xmax_cap24 VGND VPWR _0683_ net24 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_50_clk VGND VPWR clknet_3_4__leaf_clk clknet_leaf_50_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.i_regbuf\[9\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[9\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[13\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4720_ VPWR VGND VPWR VGND _1556_ _0865_ _0979_ sky130_fd_sc_hd__or2_2
XFILLER_0_17_708 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_41_clk VGND VPWR clknet_3_5__leaf_clk clknet_leaf_41_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.i_regbuf\[7\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[7\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[11\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4651_ VPWR VGND VGND VPWR _1420_ _1487_ _1486_ sky130_fd_sc_hd__nand2_1
X_7370_ VPWR VGND _3627_ i_tinyqv.cpu.instr_write_offset\[3\] _0884_ i_tinyqv.cpu.instr_data_start\[4\]
+ _3010_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_4582_ VPWR VGND VGND VPWR _1418_ i_tinyqv.cpu.instr_data\[3\]\[0\] _1417_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_6321_ VGND VPWR _2771_ _0868_ i_tinyqv.mem.qspi_data_byte_idx\[1\] i_tinyqv.mem.q_ctrl.data_ready
+ VPWR VGND sky130_fd_sc_hd__and3_1
X_6252_ VGND VPWR VPWR VGND _2728_ _0355_ _2729_ sky130_fd_sc_hd__xor2_1
X_5203_ VPWR VGND VGND VPWR _1958_ _1954_ _1956_ sky130_fd_sc_hd__or2_1
X_6183_ VGND VPWR _0343_ _2672_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5134_ VPWR VGND VGND VPWR _1890_ _1892_ _1891_ sky130_fd_sc_hd__nand2_1
X_5065_ VGND VPWR VGND VPWR _1826_ _1785_ _1804_ _1783_ _1786_ sky130_fd_sc_hd__a211o_1
X_4016_ VPWR VGND VPWR VGND i_tinyqv.cpu.data_write_n\[1\] i_tinyqv.cpu.data_read_n\[1\]
+ _0865_ _0866_ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5967_ VGND VPWR _0256_ _2543_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_32_clk VGND VPWR clknet_3_7__leaf_clk clknet_leaf_32_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_7706_ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[21\] clknet_leaf_56_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[21\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4918_ VGND VPWR _0056_ _1704_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5898_ VGND VPWR VPWR VGND _2496_ i_spi.data\[5\] _2386_ i_debug_uart_tx.uart_tx_data\[6\]
+ sky130_fd_sc_hd__mux2_1
X_7637_ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[16\] clknet_leaf_56_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[16\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.i_regbuf\[13\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[13\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[17\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4849_ VGND VPWR _0030_ _1665_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7568_ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[11\] clknet_leaf_58_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[11\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6519_ VGND VPWR VPWR VGND _2932_ i_tinyqv.mem.q_ctrl.spi_in_buffer\[1\] _2918_ i_tinyqv.mem.q_ctrl.spi_in_buffer\[5\]
+ sky130_fd_sc_hd__mux2_1
X_7499_ VGND VPWR VPWR VGND _3737_ _3736_ _2732_ _3735_ sky130_fd_sc_hd__mux2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.i_regbuf\[6\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[6\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[10\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_23_clk VGND VPWR clknet_3_6__leaf_clk clknet_leaf_23_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.i_regbuf\[4\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[4\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[8\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6870_ VGND VPWR VGND VPWR _0464_ i_tinyqv.cpu.instr_data_start\[23\] _3037_ _3238_
+ _3205_ sky130_fd_sc_hd__o211a_1
X_5821_ VGND VPWR _2447_ net200 _2448_ _2434_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_5752_ VGND VPWR _2393_ _2394_ VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_8540_ i_tinyqv.cpu.i_core.i_cycles.register\[13\] clknet_leaf_4_clk i_tinyqv.cpu.i_core.i_cycles.reg_buf\[13\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4703_ VPWR VGND VPWR VGND i_tinyqv.mem.q_ctrl.fsm_state\[1\] i_tinyqv.mem.q_ctrl.fsm_state\[0\]
+ i_tinyqv.mem.q_ctrl.fsm_state\[2\] _1539_ sky130_fd_sc_hd__or3_1
Xclkbuf_leaf_14_clk VGND VPWR clknet_3_2__leaf_clk clknet_leaf_14_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_5683_ VPWR VGND _2343_ _2337_ i_debug_uart_tx.data_to_send\[2\] VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_71_132 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_8471_ i_tinyqv.cpu.additional_mem_ops\[0\] clknet_leaf_6_clk _0569_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_7422_ VGND VPWR VPWR VGND _0726_ _3671_ _3667_ sky130_fd_sc_hd__xor2_1
X_4634_ VGND VPWR VPWR VGND net36 i_tinyqv.cpu.instr_data\[3\]\[13\] i_tinyqv.cpu.instr_data\[1\]\[13\]
+ _1470_ sky130_fd_sc_hd__mux2_2
X_7353_ VGND VPWR _3611_ _2152_ _3615_ _1439_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_4565_ VPWR VGND VPWR VGND i_tinyqv.cpu.i_core.mip\[17\] i_tinyqv.cpu.i_core.mie\[16\]
+ i_tinyqv.cpu.i_core.mip\[16\] _1401_ i_tinyqv.cpu.i_core.mie\[17\] sky130_fd_sc_hd__a22o_1
X_6304_ VGND VPWR _2761_ _2762_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_4_Right_4 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7284_ VGND VPWR _1473_ _3555_ _3560_ _2140_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_4496_ VPWR VGND VGND VPWR _1333_ _1334_ _1335_ sky130_fd_sc_hd__nor2_1
X_6235_ VPWR VGND VGND VPWR _2708_ _2713_ _2714_ sky130_fd_sc_hd__nor2_1
X_6166_ VGND VPWR _0335_ _2663_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5117_ VPWR VGND _1876_ _1875_ _1874_ VPWR VGND sky130_fd_sc_hd__and2_1
X_6097_ VGND VPWR _0313_ _2616_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5048_ VPWR VGND VGND VPWR _1806_ _1809_ _1807_ sky130_fd_sc_hd__nand2_1
X_6999_ VPWR VGND _3319_ _3318_ VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_0_23_508 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.i_regbuf\[13\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[13\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[17\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4350_ VGND VPWR VPWR VGND _1194_ gpio_out\[5\] gpio_out_sel\[5\] _1193_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_585 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4281_ VGND VPWR VPWR VGND _1128_ _1127_ _1088_ _1126_ sky130_fd_sc_hd__mux2_1
X_6020_ VGND VPWR VPWR VGND _2576_ i_tinyqv.cpu.instr_data\[2\]\[14\] _2562_ _1720_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_3_clk VGND VPWR clknet_3_0__leaf_clk clknet_leaf_3_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_7971_ i_tinyqv.cpu.i_core.cmp clknet_leaf_50_clk i_tinyqv.cpu.i_core.cmp_out VPWR
+ VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6922_ VGND VPWR VPWR VGND _0484_ _3269_ _3265_ _0691_ _3270_ net131 sky130_fd_sc_hd__a32o_1
X_6853_ VGND VPWR VPWR VGND _3223_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[30\]
+ net31 _1335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_9_513 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_5804_ VGND VPWR _0932_ _2432_ _0936_ _2433_ _0974_ _0920_ VPWR VGND sky130_fd_sc_hd__a41o_1
X_6784_ VGND VPWR VPWR VGND _3161_ _3160_ _2987_ _1590_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_313 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_3996_ VGND VPWR VGND VPWR _0847_ i_tinyqv.cpu.alu_op\[1\] _0843_ _0845_ _0846_ sky130_fd_sc_hd__a211o_2
X_5735_ _0189_ _2367_ _2371_ _2378_ _2379_ _2221_ VPWR VGND VGND VPWR sky130_fd_sc_hd__o311a_1
X_8523_ i_tinyqv.cpu.i_core.i_instrret.register\[29\] clknet_leaf_48_clk i_tinyqv.cpu.i_core.i_instrret.reg_buf\[29\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5666_ VGND VPWR _0172_ _2327_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8454_ i_tinyqv.cpu.alu_op\[0\] clknet_leaf_6_clk _0552_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_7405_ VPWR VGND VPWR VGND _3651_ _0882_ _3010_ _3657_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_349 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4617_ VGND VPWR VPWR VGND _1453_ i_tinyqv.cpu.instr_data\[3\]\[6\] _1414_ i_tinyqv.cpu.instr_data\[1\]\[6\]
+ sky130_fd_sc_hd__mux2_1
X_5597_ VGND VPWR _0151_ _2279_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8385_ i_tinyqv.cpu.data_out\[10\] clknet_leaf_26_clk _0483_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_4548_ VPWR VGND VPWR VGND _1384_ net7 sky130_fd_sc_hd__inv_2
X_7336_ VGND VPWR VGND VPWR _3603_ _3602_ _3556_ _3514_ sky130_fd_sc_hd__a21bo_1
X_4479_ VGND VPWR _1317_ _1318_ _1308_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_7267_ VPWR VGND VPWR VGND _3337_ _2121_ _3545_ _3531_ _3544_ _3546_ sky130_fd_sc_hd__a221o_2
X_6218_ VPWR VGND VPWR VGND _2026_ _2695_ _2697_ _2698_ sky130_fd_sc_hd__a21o_1
X_7198_ VPWR VGND VPWR VGND _3438_ net213 _3494_ _0536_ sky130_fd_sc_hd__a21o_1
X_6149_ VGND VPWR VPWR VGND _2654_ _2631_ _2642_ _2653_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_79_Right_79 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_75_290 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_35_121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_23_316 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_50_168 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_3850_ VPWR VGND VPWR VGND _0702_ _0698_ sky130_fd_sc_hd__inv_2
X_3781_ _0633_ net52 _0627_ net53 net56 VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
XFILLER_0_39_482 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5520_ VPWR VGND VGND VPWR _2226_ _2225_ i_uart_tx.fsm_state\[1\] _2223_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_41_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5451_ VGND VPWR _2176_ _2177_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_4402_ VPWR VGND VPWR VGND _1167_ i_tinyqv.cpu.i_core.i_shift.a\[1\] i_tinyqv.cpu.i_core.multiplier.accum\[1\]
+ _1245_ sky130_fd_sc_hd__a21oi_1
X_8170_ i_tinyqv.cpu.instr_data\[1\]\[5\] clknet_leaf_10_clk _0282_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5382_ VPWR VGND VGND VPWR _2114_ _2107_ _2113_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4333_ VGND VPWR VGND VPWR _1179_ _0830_ _1177_ _1180_ _0742_ sky130_fd_sc_hd__a2bb2o_1
X_7121_ VPWR VGND VGND VPWR _3289_ _3428_ _3427_ sky130_fd_sc_hd__nand2_1
X_4264_ VGND VPWR VPWR VGND _1111_ i_tinyqv.cpu.i_core.i_shift.a\[13\] _1028_ i_tinyqv.cpu.i_core.i_shift.a\[18\]
+ sky130_fd_sc_hd__mux2_1
X_7052_ VPWR VGND VGND VPWR _1504_ _3365_ _1461_ sky130_fd_sc_hd__nand2_1
X_6003_ VGND VPWR _0268_ _2567_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_99 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_19_Left_100 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4195_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.b\[2\] _1042_ _1041_ sky130_fd_sc_hd__nand2_1
X_7954_ i_tinyqv.cpu.i_core.time_hi\[0\] clknet_leaf_51_clk _0092_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_6905_ VPWR VGND VGND VPWR _3260_ _3261_ _2640_ sky130_fd_sc_hd__nor2_2
XFILLER_0_77_544 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_7885_ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[8\] clknet_leaf_49_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[8\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6836_ VPWR VGND VGND VPWR i_tinyqv.cpu.instr_data_start\[20\] i_tinyqv.cpu.imm\[20\]
+ _3208_ sky130_fd_sc_hd__nor2_1
X_6767_ VPWR VGND _3145_ _2995_ _1338_ VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_9_376 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_5718_ VGND VPWR _0185_ _2366_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8506_ i_tinyqv.cpu.i_core.i_instrret.register\[12\] clknet_leaf_49_clk i_tinyqv.cpu.i_core.i_instrret.reg_buf\[12\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_3979_ VGND VPWR _0779_ _0831_ _0763_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_6698_ VPWR VGND VGND VPWR _3074_ _3082_ _3037_ i_tinyqv.cpu.instr_data_start\[7\]
+ _0448_ _1753_ sky130_fd_sc_hd__o221a_1
XFILLER_0_17_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5649_ VGND VPWR _0165_ _2317_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8437_ i_tinyqv.cpu.imm\[15\] clknet_leaf_8_clk _0535_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.i_regbuf\[31\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[31\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[3\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_8368_ i_tinyqv.cpu.data_write_n\[0\] clknet_leaf_21_clk _0467_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_32_168 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold250 net279 i_tinyqv.mem.qspi_data_buf\[24\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 net290 i_tinyqv.mem.qspi_data_buf\[30\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_7319_ VGND VPWR VPWR VGND _3589_ _0662_ _2153_ _3588_ sky130_fd_sc_hd__mux2_1
X_8299_ i_tinyqv.mem.q_ctrl.nibbles_remaining\[2\] clknet_leaf_14_clk _0398_ VPWR
+ VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold272 net301 i_tinyqv.mem.q_ctrl.addr\[17\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 net312 i_tinyqv.mem.q_ctrl.addr\[8\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.i_regbuf\[27\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[27\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[31\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.i_regbuf\[16\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[16\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[20\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_422 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_24_614 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_36_485 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_instrret.i_regbuf\[26\] i_tinyqv.cpu.i_core.i_instrret.reg_buf\[26\]
+ i_tinyqv.cpu.i_core.i_instrret.register\[30\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xinput7 VPWR VGND VPWR VGND net7 ui_in[5] sky130_fd_sc_hd__dlymetal6s2s_1
X_4951_ VGND VPWR _1731_ gpio_out\[0\] _1729_ _1730_ VPWR VGND sky130_fd_sc_hd__and3_1
X_3902_ VPWR VGND VPWR VGND _0613_ i_tinyqv.cpu.instr_data_start\[17\] _0753_ _0754_
+ sky130_fd_sc_hd__a21oi_1
X_7670_ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[17\] clknet_leaf_55_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[17\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4882_ VGND VPWR VPWR VGND _1684_ i_tinyqv.cpu.debug_rd\[3\] _1680_ i_tinyqv.cpu.i_core.i_registers.reg_access\[7\]\[3\]
+ sky130_fd_sc_hd__mux2_1
X_6621_ VGND VPWR VPWR VGND _3015_ _3014_ _3012_ i_tinyqv.cpu.data_addr\[2\] sky130_fd_sc_hd__mux2_1
X_3833_ VPWR VGND VPWR VGND _0684_ i_tinyqv.cpu.i_core.i_registers.reg_access\[1\]\[3\]
+ net24 _0685_ i_tinyqv.cpu.i_core.i_registers.reg_access\[13\]\[3\] sky130_fd_sc_hd__a22o_1
X_6552_ VPWR VGND VGND VPWR _2961_ i_debug_uart_tx.uart_tx_data\[5\] _2909_ sky130_fd_sc_hd__or2_1
X_3764_ VPWR VGND _0616_ i_tinyqv.cpu.counter\[2\] i_tinyqv.cpu.counter\[3\] VPWR
+ VGND sky130_fd_sc_hd__and2_1
X_6483_ VGND VPWR _0414_ _2901_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5503_ VGND VPWR _2212_ _2200_ _2214_ net157 VPWR VGND sky130_fd_sc_hd__o21ai_1
X_8222_ i_tinyqv.cpu.i_core.multiplier.accum\[5\] clknet_leaf_44_clk _0023_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5434_ _2162_ _2160_ _1752_ _2152_ _2161_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
X_8153_ i_tinyqv.cpu.instr_data\[2\]\[2\] clknet_leaf_11_clk _0265_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5365_ VGND VPWR VGND VPWR net43 _2099_ _2089_ sky130_fd_sc_hd__or2b_1
X_7104_ VGND VPWR VGND VPWR _3413_ _3409_ _3410_ _3364_ _3412_ sky130_fd_sc_hd__a211o_1
X_8084_ gpio_out_sel\[3\] clknet_leaf_18_clk _0011_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5296_ VGND VPWR i_tinyqv.cpu.i_core.cy_out _2046_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4316_ VPWR VGND _1163_ _1162_ _1144_ _1046_ _1121_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_4247_ VGND VPWR VPWR VGND _1094_ i_tinyqv.cpu.i_core.i_shift.a\[25\] _1036_ i_tinyqv.cpu.i_core.i_shift.a\[6\]
+ sky130_fd_sc_hd__mux2_1
X_7035_ VPWR VGND VGND VPWR _1468_ _3297_ _3349_ sky130_fd_sc_hd__nor2_1
X_4178_ VPWR VGND VGND VPWR _0852_ _1025_ _0849_ sky130_fd_sc_hd__nand2_1
X_7937_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[28\] clknet_leaf_49_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[28\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7868_ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[23\] clknet_leaf_47_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[23\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6819_ VPWR VGND VPWR VGND _3185_ _3039_ _3193_ _2306_ _1345_ _3192_ sky130_fd_sc_hd__a221o_1
X_7799_ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[18\] clknet_leaf_57_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[18\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.i_regbuf\[28\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[28\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.i_regbuf\[17\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[17\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[21\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_56_525 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_71_528 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.i_regbuf\[31\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[31\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[3\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_411 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_5150_ VPWR VGND VGND VPWR _1905_ _1907_ _1906_ sky130_fd_sc_hd__nand2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.i_regbuf\[20\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[20\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[24\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5081_ VGND VPWR _1840_ _1841_ i_tinyqv.cpu.i_core.multiplier.accum\[7\] VPWR VGND
+ sky130_fd_sc_hd__xnor2_1
X_4101_ VPWR VGND VGND VPWR _0922_ _0937_ _0840_ _0948_ sky130_fd_sc_hd__nor3_1
X_4032_ VPWR VGND _0879_ i_tinyqv.cpu.is_lui _0653_ VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_2_56 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_5983_ VGND VPWR _0261_ _2554_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4934_ VGND VPWR VGND VPWR _1709_ i_tinyqv.mem.q_ctrl.nibbles_remaining\[0\] _1715_
+ _1718_ i_tinyqv.mem.q_ctrl.addr\[21\] sky130_fd_sc_hd__a2bb2o_1
X_7722_ i_tinyqv.cpu.i_core.i_registers.reg_access\[9\]\[1\] clknet_leaf_54_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[5\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XANTENNA_23 i_tinyqv.mem.q_ctrl.addr\[21\] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_12 i_tinyqv.cpu.i_core.imm_lo\[5\] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_7653_ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[0\] clknet_leaf_56_clk _0038_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4865_ VGND VPWR VGND VPWR _1674_ _1658_ _1640_ i_tinyqv.cpu.i_core.i_registers.rd\[1\]
+ sky130_fd_sc_hd__and3b_2
XFILLER_0_74_399 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4796_ VGND VPWR VGND VPWR i_tinyqv.mem.qspi_data_buf\[31\] i_tinyqv.mem.qspi_data_buf\[27\]
+ _0974_ i_tinyqv.cpu.instr_data_in\[15\] i_tinyqv.cpu.instr_data_in\[11\] _0979_
+ _1631_ sky130_fd_sc_hd__mux4_1
X_6604_ VGND VPWR VPWR VGND _3001_ _3000_ _2991_ _2507_ sky130_fd_sc_hd__mux2_1
XANTENNA_45 i_tinyqv.cpu.i_core.imm_lo\[9\] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_7584_ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[27\] clknet_leaf_59_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[27\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_3816_ VPWR VGND VGND VPWR _0662_ _0663_ _0660_ i_tinyqv.cpu.i_core.i_registers.rs2\[3\]
+ _0668_ sky130_fd_sc_hd__and4b_2
XANTENNA_34 i_tinyqv.cpu.i_core.imm_lo\[9\] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_6535_ VGND VPWR VPWR VGND _2946_ _2945_ _2929_ _2944_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_499 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6466_ VPWR VGND VGND VPWR _1181_ _2625_ _2890_ sky130_fd_sc_hd__nor2_1
X_8205_ i_tinyqv.cpu.i_core.i_shift.a\[24\] clknet_leaf_40_clk _0317_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_6397_ VGND VPWR _2835_ _2833_ _2832_ _2834_ VPWR VGND sky130_fd_sc_hd__and3_1
X_5417_ VGND VPWR _2146_ _2147_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_5348_ VGND VPWR VPWR VGND _2086_ i_tinyqv.cpu.i_core.interrupt_req\[1\] _2084_ i_tinyqv.cpu.i_core.last_interrupt_req\[1\]
+ sky130_fd_sc_hd__mux2_1
X_8136_ i_tinyqv.cpu.data_addr\[11\] clknet_leaf_33_clk _0248_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_8067_ i_spi.read_latency clknet_leaf_27_clk _0202_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5279_ VGND VPWR VPWR VGND _2028_ _2031_ _2030_ sky130_fd_sc_hd__xor2_1
X_7018_ VPWR VGND VGND VPWR _3334_ _3319_ _3335_ sky130_fd_sc_hd__nor2_1
Xmax_cap14 VPWR VGND net14 _1003_ VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_0_80_358 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_61_561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.i_regbuf\[9\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[9\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[13\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4650_ VGND VPWR VPWR VGND _1486_ _1408_ _1485_ _1484_ sky130_fd_sc_hd__mux2_4
Xinput10 VGND VPWR net10 uio_in[1] VPWR VGND sky130_fd_sc_hd__buf_1
X_6320_ VGND VPWR _0382_ _2770_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4581_ VGND VPWR _1411_ _1410_ _1417_ net325 VPWR VGND sky130_fd_sc_hd__o21ai_2
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.i_regbuf\[21\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[21\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[25\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6251_ _2729_ _2708_ _2713_ _2722_ _2723_ VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_5202_ VPWR VGND VGND VPWR _1954_ _1957_ _1956_ sky130_fd_sc_hd__nand2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.i_regbuf\[7\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[7\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[11\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6182_ VGND VPWR VPWR VGND _2672_ i_tinyqv.cpu.i_core.mepc\[18\] _2667_ i_tinyqv.cpu.i_core.mepc\[14\]
+ sky130_fd_sc_hd__mux2_1
X_5133_ VPWR VGND VGND VPWR _1877_ _1862_ _1891_ _1889_ sky130_fd_sc_hd__nand3_1
X_5064_ VGND VPWR _1824_ _1825_ _1822_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_4015_ VPWR VGND VPWR VGND i_tinyqv.cpu.data_addr\[26\] i_tinyqv.cpu.data_addr\[25\]
+ i_tinyqv.cpu.data_addr\[27\] _0865_ sky130_fd_sc_hd__or3_4
X_5966_ VGND VPWR VPWR VGND _2543_ _2542_ _2524_ i_tinyqv.cpu.data_addr\[19\] sky130_fd_sc_hd__mux2_1
X_5897_ VGND VPWR _0234_ _2495_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7705_ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[20\] clknet_leaf_0_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[20\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4917_ VGND VPWR VPWR VGND _1704_ _1380_ _1701_ i_tinyqv.cpu.i_core.i_registers.reg_access\[1\]\[2\]
+ sky130_fd_sc_hd__mux2_1
X_7636_ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[15\] clknet_leaf_45_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[15\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4848_ VGND VPWR VPWR VGND _1665_ i_tinyqv.cpu.debug_rd\[0\] _1664_ i_tinyqv.cpu.i_core.i_registers.reg_access\[10\]\[0\]
+ sky130_fd_sc_hd__mux2_1
X_7567_ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[10\] clknet_leaf_54_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[10\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4779_ VPWR VGND VPWR VGND _1603_ _0697_ _0880_ _1614_ _1613_ sky130_fd_sc_hd__a22o_1
X_6518_ VGND VPWR VPWR VGND _2931_ _2930_ _2916_ net11 sky130_fd_sc_hd__mux2_1
X_7498_ VGND VPWR VPWR VGND _3736_ i_tinyqv.mem.q_ctrl.addr\[19\] _3007_ i_tinyqv.mem.q_ctrl.addr\[23\]
+ sky130_fd_sc_hd__mux2_1
X_6449_ VPWR VGND _2878_ _2877_ VPWR VGND sky130_fd_sc_hd__buf_4
X_8119_ i_spi.data\[2\] clknet_leaf_19_clk _0231_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.i_regbuf\[6\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[6\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[10\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_572 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_34_583 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_21_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_29_300 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5820_ _2447_ net42 _2088_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_5751_ i_spi.busy _1000_ _2393_ _1557_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_4702_ VGND VPWR VGND VPWR _1538_ i_tinyqv.mem.q_ctrl.data_ready i_tinyqv.mem.q_ctrl.data_req
+ _1385_ _0872_ sky130_fd_sc_hd__o211a_1
X_8470_ i_tinyqv.cpu.instr_len\[2\] clknet_leaf_7_clk _0568_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5682_ VGND VPWR VGND VPWR _0173_ net117 _2330_ _2342_ _2299_ sky130_fd_sc_hd__o211a_1
X_7421_ VPWR VGND VPWR VGND net302 _3007_ _0583_ _3009_ net303 _3670_ sky130_fd_sc_hd__a221o_1
X_4633_ VPWR VGND VGND VPWR _1469_ _1420_ _1468_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_358 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_4564_ VGND VPWR VPWR VGND i_tinyqv.cpu.i_core.i_cycles.rstn _1400_ sky130_fd_sc_hd__clkinv_4
X_7352_ VGND VPWR VGND VPWR _0570_ net242 _2152_ _3614_ _1753_ sky130_fd_sc_hd__o211a_1
X_6303_ _0868_ i_tinyqv.mem.q_ctrl.data_ready _2761_ i_tinyqv.mem.qspi_data_byte_idx\[1\]
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_7283_ VGND VPWR _0556_ _3559_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6234_ VGND VPWR VPWR VGND _2710_ _2711_ _2713_ _2041_ sky130_fd_sc_hd__a21boi_2
X_4495_ VPWR VGND VPWR VGND _0900_ i_tinyqv.cpu.instr_data_start\[21\] i_tinyqv.cpu.instr_data_start\[22\]
+ _1334_ sky130_fd_sc_hd__a21oi_1
X_6165_ VGND VPWR VPWR VGND _2663_ i_tinyqv.cpu.i_core.mepc\[10\] _2656_ i_tinyqv.cpu.i_core.mepc\[6\]
+ sky130_fd_sc_hd__mux2_1
X_5116_ VPWR VGND VPWR VGND _1851_ _1873_ _1853_ _1875_ sky130_fd_sc_hd__or3_1
X_6096_ VGND VPWR VPWR VGND _2616_ i_tinyqv.cpu.i_core.i_shift.a\[20\] _2595_ i_tinyqv.cpu.i_core.i_shift.a\[24\]
+ sky130_fd_sc_hd__mux2_1
X_5047_ VPWR VGND VGND VPWR _1808_ _1806_ _1807_ sky130_fd_sc_hd__or2_1
X_6998_ VGND VPWR VPWR VGND _1492_ _1452_ _1491_ _3318_ sky130_fd_sc_hd__or3b_1
X_5949_ VGND VPWR _0250_ _2531_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_163 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_62_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_7619_ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[30\] clknet_leaf_2_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[30\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.i_regbuf\[21\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[21\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[25\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.i_regbuf\[10\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[10\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[14\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4280_ VGND VPWR VPWR VGND _1127_ _1071_ _1103_ _1069_ sky130_fd_sc_hd__mux2_1
X_7970_ i_tinyqv.cpu.i_core.i_registers.rd\[3\] clknet_leaf_6_clk _0107_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_6921_ VGND VPWR VPWR VGND _0483_ _3268_ _3265_ _0691_ _3270_ net132 sky130_fd_sc_hd__a32o_1
X_6852_ VGND VPWR VGND VPWR _0462_ i_tinyqv.cpu.instr_data_start\[21\] _3123_ _3222_
+ _3205_ sky130_fd_sc_hd__o211a_1
X_5803_ VPWR VGND VPWR VGND _2432_ _0942_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_461 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_6783_ VPWR VGND VPWR VGND _3160_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[23\]
+ sky130_fd_sc_hd__inv_2
X_8522_ i_tinyqv.cpu.i_core.i_instrret.register\[28\] clknet_leaf_49_clk i_tinyqv.cpu.i_core.i_instrret.reg_buf\[28\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_3995_ VPWR VGND i_tinyqv.cpu.alu_op\[1\] _0846_ i_tinyqv.cpu.alu_op\[3\] VPWR VGND
+ sky130_fd_sc_hd__and2_2
XFILLER_0_45_612 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5734_ VPWR VGND VGND VPWR _2379_ i_debug_uart_tx.fsm_state\[3\] _2375_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_122 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5665_ VGND VPWR VPWR VGND _2327_ _1721_ _2308_ net281 sky130_fd_sc_hd__mux2_1
X_8453_ i_tinyqv.cpu.imm\[31\] clknet_leaf_22_clk _0551_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_369 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_8384_ i_spi.dc_in clknet_leaf_26_clk _0482_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7404_ VPWR VGND VGND VPWR _3656_ _0882_ _3651_ sky130_fd_sc_hd__or2_1
X_4616_ VGND VPWR VPWR VGND _1409_ _1451_ _1450_ _1452_ sky130_fd_sc_hd__mux2_2
X_5596_ VPWR VGND VGND VPWR _2279_ _2229_ _2239_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_7335_ VGND VPWR VGND VPWR _3602_ _2125_ _1487_ _1426_ _3304_ sky130_fd_sc_hd__a211o_1
X_4547_ VGND VPWR _1383_ uo_out[3] VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_4478_ VGND VPWR _1316_ _1317_ i_tinyqv.cpu.i_core.multiplier.accum\[2\] VPWR VGND
+ sky130_fd_sc_hd__xnor2_1
X_7266_ VPWR VGND VGND VPWR _3545_ _3304_ _3539_ sky130_fd_sc_hd__or2_1
X_6217_ VGND VPWR _2696_ _2697_ _2694_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_7197_ VGND VPWR _3494_ _3492_ _3359_ _3493_ VPWR VGND sky130_fd_sc_hd__and3_1
X_6148_ VPWR VGND VGND VPWR _0956_ _0693_ _0696_ _2653_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_13_Left_94 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6079_ VGND VPWR _0304_ _2607_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_206 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_3780_ VGND VPWR VGND VPWR _0631_ _0629_ _0630_ _0632_ i_tinyqv.cpu.i_core.i_registers.reg_access\[12\]\[3\]
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_39_494 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5450_ VGND VPWR _2176_ _2170_ _0990_ _2175_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_2_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_4401_ VGND VPWR _1244_ i_tinyqv.cpu.i_core.multiplier.accum\[1\] i_tinyqv.cpu.i_core.i_shift.a\[1\]
+ _1166_ VPWR VGND sky130_fd_sc_hd__and3_1
X_5381_ VGND VPWR VPWR VGND _2113_ i_tinyqv.cpu.i_core.mstatus_mie _2112_ _2103_ sky130_fd_sc_hd__mux2_1
X_4332_ VPWR VGND VGND VPWR _0708_ net79 _1178_ _1179_ sky130_fd_sc_hd__o21a_1
X_7120_ VPWR VGND VGND VPWR _3367_ i_tinyqv.cpu.instr_data\[1\]\[10\] _3365_ i_tinyqv.cpu.instr_data\[0\]\[10\]
+ _3427_ _3426_ sky130_fd_sc_hd__o221a_1
X_4263_ VGND VPWR VPWR VGND _1110_ i_tinyqv.cpu.i_core.i_shift.a\[12\] _1028_ i_tinyqv.cpu.i_core.i_shift.a\[19\]
+ sky130_fd_sc_hd__mux2_1
X_7051_ VPWR VGND _3364_ _3363_ VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_0_10_589 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_6002_ VGND VPWR VPWR VGND _2567_ i_tinyqv.cpu.instr_data\[2\]\[5\] _2563_ i_tinyqv.cpu.instr_data_in\[5\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_64 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4194_ VGND VPWR _1027_ _1041_ _0838_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_7953_ i_tinyqv.cpu.i_core.is_double_fault_r clknet_leaf_37_clk _0091_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6904_ VPWR VGND VGND VPWR _3260_ _1026_ _0955_ sky130_fd_sc_hd__nand2_2
XFILLER_0_77_556 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7884_ i_tinyqv.cpu.i_core.i_registers.reg_access\[2\]\[3\] clknet_leaf_48_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[7\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6835_ VPWR VGND VPWR VGND _3195_ _3207_ _3196_ _3198_ sky130_fd_sc_hd__a21boi_1
X_6766_ VGND VPWR VGND VPWR _0454_ i_tinyqv.cpu.instr_data_start\[13\] _3123_ _3144_
+ _3093_ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_355 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_3978_ VGND VPWR VPWR VGND _0742_ _0830_ _0829_ sky130_fd_sc_hd__xor2_1
X_5717_ VGND VPWR _2366_ _1729_ i_debug_uart_tx.cycle_counter\[4\] _2364_ VPWR VGND
+ sky130_fd_sc_hd__and3_1
X_8505_ i_tinyqv.cpu.i_core.i_instrret.register\[11\] clknet_leaf_45_clk i_tinyqv.cpu.i_core.i_instrret.reg_buf\[11\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_656 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6697_ VPWR VGND _3082_ _3081_ _3075_ _3051_ _3028_ VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_18_689 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_8436_ i_tinyqv.cpu.imm\[14\] clknet_leaf_21_clk _0534_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_5648_ VGND VPWR VPWR VGND _2317_ _2316_ _2309_ i_tinyqv.cpu.instr_data\[3\]\[8\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_561 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_32_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5579_ VPWR VGND VGND VPWR _2268_ i_uart_rx.recieved_data\[3\] _2264_ sky130_fd_sc_hd__or2_1
X_8367_ i_tinyqv.cpu.was_early_branch clknet_leaf_24_clk _0466_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_2
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.i_regbuf\[24\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[24\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[28\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_8298_ i_tinyqv.mem.q_ctrl.nibbles_remaining\[1\] clknet_leaf_14_clk _0397_ VPWR
+ VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold240 net269 i_tinyqv.mem.data_from_read\[18\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 net280 i_tinyqv.mem.data_from_read\[16\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 net291 i_tinyqv.cpu.instr_data\[0\]\[3\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7318_ VPWR VGND VGND VPWR _2147_ _3585_ _3587_ _3588_ sky130_fd_sc_hd__o21a_1
Xhold284 net313 i_debug_uart_tx.uart_tx_data\[5\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 net302 i_tinyqv.mem.q_ctrl.addr\[7\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7249_ VPWR VGND VGND VPWR _2140_ _1466_ _3530_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_464 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_23_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xinput8 VGND VPWR net8 ui_in[6] VPWR VGND sky130_fd_sc_hd__buf_1
Xi_tinyqv.cpu.i_core.i_instrret.i_regbuf\[19\] i_tinyqv.cpu.i_core.i_instrret.reg_buf\[19\]
+ i_tinyqv.cpu.i_core.i_instrret.register\[23\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_512 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_4950_ VPWR VGND VGND VPWR _1730_ _1001_ _1725_ sky130_fd_sc_hd__nand2_2
X_3901_ VPWR VGND VPWR VGND _0751_ i_tinyqv.cpu.instr_data_start\[21\] _0610_ _0753_
+ _0752_ sky130_fd_sc_hd__a22o_1
X_4881_ VGND VPWR _0072_ _1683_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6620_ VGND VPWR VPWR VGND _3014_ _3000_ _3010_ i_tinyqv.cpu.instr_write_offset\[2\]
+ sky130_fd_sc_hd__mux2_1
X_3832_ VPWR VGND VGND VPWR _0663_ _0660_ _0661_ _0662_ _0684_ sky130_fd_sc_hd__and4b_2
X_6551_ VGND VPWR VPWR VGND _2960_ i_tinyqv.cpu.data_out\[21\] _2912_ i_tinyqv.cpu.data_out\[29\]
+ sky130_fd_sc_hd__mux2_1
X_5502_ VPWR VGND VGND VPWR _2212_ _2213_ _0122_ sky130_fd_sc_hd__nor2_1
X_3763_ VPWR VGND VGND VPWR _0608_ _0615_ _0614_ sky130_fd_sc_hd__nor2_2
X_6482_ VGND VPWR VPWR VGND _2901_ i_tinyqv.mem.q_ctrl.spi_in_buffer\[3\] _2897_ net13
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_136 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_8221_ i_tinyqv.cpu.i_core.multiplier.accum\[4\] clknet_leaf_45_clk _0022_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5433_ VPWR VGND VPWR VGND _1501_ _2137_ _2161_ _2141_ _1491_ _2149_ sky130_fd_sc_hd__a221o_1
X_8152_ i_tinyqv.cpu.data_addr\[27\] clknet_leaf_35_clk _0264_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_5364_ VPWR VGND VPWR VGND _2087_ net223 _0840_ _0099_ _2098_ sky130_fd_sc_hd__a22o_1
X_4315_ VGND VPWR VGND VPWR _1048_ _1161_ _1077_ _1148_ _1153_ _1162_ sky130_fd_sc_hd__a311o_1
X_7103_ VPWR VGND VPWR VGND _3412_ _2121_ _2130_ _3411_ _3305_ _3377_ sky130_fd_sc_hd__o32a_1
X_8083_ gpio_out_sel\[2\] clknet_leaf_18_clk _0010_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5295_ VPWR VGND _2046_ _0821_ _0701_ VPWR VGND sky130_fd_sc_hd__and2_1
X_4246_ VGND VPWR VPWR VGND _1093_ i_tinyqv.cpu.i_core.i_shift.a\[24\] _1036_ _1054_
+ sky130_fd_sc_hd__mux2_1
X_7034_ VPWR VGND VGND VPWR _3346_ _3348_ _3347_ sky130_fd_sc_hd__nand2_1
X_4177_ VPWR VGND VPWR VGND _1021_ _0955_ _1023_ _1024_ sky130_fd_sc_hd__a21o_1
X_7936_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[27\] clknet_leaf_36_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[27\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7867_ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[22\] clknet_leaf_3_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[22\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6818_ VGND VPWR VGND VPWR _3192_ _3040_ _3190_ _3191_ net40 sky130_fd_sc_hd__o211a_1
X_7798_ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[17\] clknet_leaf_1_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[17\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6749_ VGND VPWR _3128_ _3129_ _3125_ VPWR VGND sky130_fd_sc_hd__xnor2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.i_regbuf\[25\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[25\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[29\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_8419_ i_tinyqv.cpu.is_jalr clknet_leaf_7_clk _0517_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_38_Left_119 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_52_710 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.i_regbuf\[24\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[24\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[28\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_47_Left_128 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_cycles.i_regbuf\[22\] i_tinyqv.cpu.i_core.i_cycles.reg_buf\[22\]
+ i_tinyqv.cpu.i_core.i_cycles.register\[26\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_684 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_5080_ VPWR VGND _1840_ _1839_ _1838_ VPWR VGND sky130_fd_sc_hd__and2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.i_regbuf\[13\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[13\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[17\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4100_ VPWR VGND VGND VPWR _0937_ _0928_ _0946_ _0947_ sky130_fd_sc_hd__nor3_1
X_4031_ VPWR VGND VGND VPWR _0878_ i_tinyqv.cpu.data_ready_core _0851_ sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_56_Left_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5982_ VPWR VGND _2554_ _2553_ _2079_ VPWR VGND sky130_fd_sc_hd__and2_1
X_4933_ VPWR VGND _1717_ i_tinyqv.cpu.instr_data_in\[13\] VPWR VGND sky130_fd_sc_hd__buf_2
X_7721_ i_tinyqv.cpu.i_core.i_registers.reg_access\[9\]\[0\] clknet_leaf_1_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[4\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4864_ VGND VPWR _0081_ _1673_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7652_ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[31\] clknet_leaf_46_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[31\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XANTENNA_13 i_tinyqv.cpu.i_core.imm_lo\[9\] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_24 i_uart_rx.recieved_data\[7\] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_4795_ VPWR VGND _1630_ _1629_ _1626_ _0689_ _0956_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_6603_ VPWR VGND VGND VPWR _2998_ _2999_ _3000_ sky130_fd_sc_hd__nor2_1
XANTENNA_46 i_tinyqv.cpu.i_core.imm_lo\[9\] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_35 i_tinyqv.cpu.i_core.imm_lo\[9\] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_7583_ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[26\] clknet_leaf_55_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[26\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_3815_ VPWR VGND VGND VPWR _0667_ net39 _0663_ sky130_fd_sc_hd__nor2b_2
X_6534_ VGND VPWR VPWR VGND _2945_ i_tinyqv.cpu.data_out\[11\] _2909_ i_debug_uart_tx.uart_tx_data\[3\]
+ sky130_fd_sc_hd__mux2_1
X_6465_ VPWR VGND VPWR VGND _2888_ _1540_ _2889_ _0408_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_65_Left_146 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_70_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_8204_ i_tinyqv.cpu.i_core.i_shift.a\[23\] clknet_leaf_40_clk _0316_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5416_ VGND VPWR VGND VPWR _1439_ _2146_ _1440_ sky130_fd_sc_hd__or2b_1
X_6396_ VGND VPWR _2834_ _1711_ _1713_ _2794_ VPWR VGND sky130_fd_sc_hd__and3_1
X_5347_ VGND VPWR _0095_ net251 VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8135_ i_tinyqv.cpu.data_addr\[10\] clknet_leaf_34_clk _0247_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_11_662 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_8066_ i_debug_uart_tx.txd_reg clknet_leaf_30_clk _0201_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5278_ VGND VPWR _2001_ _2029_ _2030_ _2000_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_4229_ VPWR VGND VPWR VGND _1045_ _1038_ _1044_ _1076_ sky130_fd_sc_hd__a21o_1
X_7017_ VPWR VGND VPWR VGND _3334_ _1455_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_74_Left_155 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xmax_cap26 VGND VPWR net26 _0638_ VPWR VGND sky130_fd_sc_hd__buf_1
Xmax_cap15 VGND VPWR net15 _0943_ VPWR VGND sky130_fd_sc_hd__buf_1
X_7919_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[10\] clknet_leaf_26_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[10\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_710 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_46_592 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_61_540 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_0_309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_1_Left_82 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xinput11 VGND VPWR net11 uio_in[2] VPWR VGND sky130_fd_sc_hd__buf_1
X_4580_ VGND VPWR VPWR VGND _1416_ _0653_ _1415_ _0749_ sky130_fd_sc_hd__mux2_4
XFILLER_0_52_540 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_4_626 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_24_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_3_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6250_ VGND VPWR _2727_ _2728_ _2725_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_5201_ VGND VPWR _1927_ _1955_ _1956_ _1926_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_6181_ VGND VPWR _0342_ _2671_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.i_regbuf\[14\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[14\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[18\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5132_ VPWR VGND VPWR VGND _1862_ _1877_ _1889_ _1890_ sky130_fd_sc_hd__a21o_1
X_5063_ VGND VPWR VGND VPWR _1823_ _1800_ _1801_ _1824_ sky130_fd_sc_hd__o21ba_1
X_4014_ VPWR VGND VPWR VGND _0864_ i_tinyqv.mem.qspi_data_byte_idx\[1\] sky130_fd_sc_hd__inv_2
X_5965_ VGND VPWR VPWR VGND _2542_ i_tinyqv.cpu.i_core.mepc\[19\] _2107_ i_tinyqv.cpu.i_core.i_shift.a\[23\]
+ sky130_fd_sc_hd__mux2_1
X_5896_ VGND VPWR VPWR VGND _2495_ _2494_ _2399_ i_spi.data\[5\] sky130_fd_sc_hd__mux2_1
X_7704_ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[19\] clknet_leaf_58_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[19\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4916_ VGND VPWR _0055_ _1703_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7635_ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[14\] clknet_leaf_45_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[14\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4847_ VPWR VGND _1641_ _1664_ _1658_ VPWR VGND sky130_fd_sc_hd__and2_2
X_7566_ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[9\] clknet_leaf_58_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[9\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4778_ VPWR VGND VPWR VGND _1612_ _0921_ _0880_ _1613_ sky130_fd_sc_hd__a21oi_1
X_6517_ VGND VPWR VPWR VGND _2930_ _2928_ _2929_ _2927_ sky130_fd_sc_hd__mux2_1
X_7497_ VGND VPWR VPWR VGND _3735_ _3734_ _2681_ i_tinyqv.cpu.data_addr\[23\] sky130_fd_sc_hd__mux2_1
XFILLER_0_43_595 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6448_ VGND VPWR _2734_ _2877_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xi_tinyqv.cpu.i_core.i_instrret.i_regbuf\[8\] i_tinyqv.cpu.i_core.i_instrret.reg_buf\[8\]
+ i_tinyqv.cpu.i_core.i_instrret.register\[12\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6379_ VGND VPWR VPWR VGND _2819_ _2818_ _2804_ _2815_ sky130_fd_sc_hd__mux2_1
X_8118_ i_spi.data\[1\] clknet_leaf_27_clk _0230_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_8049_ i_debug_uart_tx.cycle_counter\[3\] clknet_leaf_30_clk _0184_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_654 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_38_378 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_1_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_5750_ VPWR VGND _2392_ _2383_ i_spi.busy VPWR VGND sky130_fd_sc_hd__and2_1
X_5681_ VGND VPWR VGND VPWR _2342_ _2336_ _2338_ i_debug_uart_tx.data_to_send\[0\]
+ _2341_ sky130_fd_sc_hd__a211o_1
X_4701_ VPWR VGND VPWR VGND _1530_ _1535_ _1536_ _1537_ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_635 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_7420_ VGND VPWR VGND VPWR _3670_ net96 _3012_ _3004_ _3669_ sky130_fd_sc_hd__o211a_1
X_4632_ VGND VPWR VGND VPWR _1425_ _1461_ _1421_ _1423_ _1468_ sky130_fd_sc_hd__a31o_2
X_4563_ VPWR VGND VGND VPWR _1398_ _1399_ sky130_fd_sc_hd__buf_8
XFILLER_0_8_45 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_7351_ VGND VPWR VGND VPWR _3614_ _3613_ _3610_ _2152_ sky130_fd_sc_hd__a21bo_1
X_6302_ VGND VPWR _0374_ _2760_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7282_ VGND VPWR VPWR VGND _3559_ _3558_ _3395_ i_tinyqv.cpu.i_core.mem_op\[0\] sky130_fd_sc_hd__mux2_1
X_4494_ VGND VPWR _1333_ i_tinyqv.cpu.instr_data_start\[21\] i_tinyqv.cpu.instr_data_start\[22\]
+ _0900_ VPWR VGND sky130_fd_sc_hd__and3_1
X_6233_ VGND VPWR VPWR VGND _2710_ _0353_ _2712_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_6164_ VGND VPWR _0334_ _2662_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5115_ VGND VPWR _1851_ _1873_ _1874_ _1853_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_6095_ VGND VPWR _0312_ _2615_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5046_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[4\] _1807_ _1309_ sky130_fd_sc_hd__nand2_1
X_6997_ VPWR VGND VGND VPWR _2067_ _3317_ _0512_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5948_ VGND VPWR VPWR VGND _2531_ _2530_ _2524_ i_tinyqv.cpu.data_addr\[13\] sky130_fd_sc_hd__mux2_1
X_5879_ VPWR VGND VPWR VGND _2484_ _2309_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_261 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7618_ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[29\] clknet_leaf_52_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[29\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.i_regbuf\[4\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[4\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[8\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_16_551 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7549_ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[24\] clknet_leaf_47_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[24\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.i_regbuf\[14\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[14\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[18\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6920_ VGND VPWR VPWR VGND _0482_ _3267_ _3265_ _0691_ _3270_ net169 sky130_fd_sc_hd__a32o_1
X_6851_ VPWR VGND VPWR VGND _3220_ _3051_ _3221_ _3222_ sky130_fd_sc_hd__a21o_1
X_5802_ VPWR VGND VPWR VGND _2431_ net192 sky130_fd_sc_hd__inv_2
X_6782_ VGND VPWR VPWR VGND _3159_ _3158_ _2991_ _2534_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_548 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_8521_ i_tinyqv.cpu.i_core.i_instrret.register\[27\] clknet_leaf_46_clk i_tinyqv.cpu.i_core.i_instrret.reg_buf\[27\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_3994_ VPWR VGND _0845_ i_tinyqv.cpu.alu_op\[0\] _0844_ VPWR VGND sky130_fd_sc_hd__and2_1
X_5733_ VGND VPWR VPWR VGND i_debug_uart_tx.fsm_state\[2\] _2378_ i_debug_uart_tx.fsm_state\[0\]
+ sky130_fd_sc_hd__xor2_1
X_5664_ VGND VPWR _0171_ _2326_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_8452_ i_tinyqv.cpu.imm\[30\] clknet_leaf_22_clk _0550_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5595_ VGND VPWR VGND VPWR _0150_ net191 _2277_ _2278_ _2182_ sky130_fd_sc_hd__o211a_1
X_8383_ i_spi.end_txn clknet_leaf_26_clk _0481_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7403_ VPWR VGND VPWR VGND _3655_ _3653_ _3654_ _0580_ _2733_ sky130_fd_sc_hd__a22o_1
X_4615_ VGND VPWR VPWR VGND _1451_ i_tinyqv.cpu.instr_data\[2\]\[5\] _1449_ i_tinyqv.cpu.instr_data\[0\]\[5\]
+ sky130_fd_sc_hd__mux2_1
X_4546_ VGND VPWR VPWR VGND _1383_ gpio_out\[3\] gpio_out_sel\[3\] _1382_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_543 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7334_ VGND VPWR VPWR VGND _0661_ _3601_ _3595_ sky130_fd_sc_hd__xor2_1
X_4477_ VPWR VGND VGND VPWR _1310_ _1314_ _1315_ _1316_ sky130_fd_sc_hd__o21a_1
X_7265_ VGND VPWR VGND VPWR _3544_ _3533_ _2124_ _3540_ sky130_fd_sc_hd__a21bo_1
X_6216_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[14\] _2696_ _1880_ sky130_fd_sc_hd__nand2_1
X_7196_ VGND VPWR VGND VPWR _3493_ _3331_ _3470_ _3305_ _3481_ sky130_fd_sc_hd__a211o_1
X_6147_ VGND VPWR _0327_ _2652_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6078_ VGND VPWR VPWR VGND _2607_ _1060_ _2593_ i_tinyqv.cpu.i_core.i_shift.a\[11\]
+ sky130_fd_sc_hd__mux2_1
X_5029_ VPWR VGND _1791_ _1789_ _1767_ i_tinyqv.cpu.i_core.i_shift.a\[3\] _1790_ VGND
+ VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_51_605 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_36_657 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_51_649 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_26_101 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_27_613 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_6_529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4400_ VPWR VGND VPWR VGND _1242_ _0955_ _1023_ _1243_ sky130_fd_sc_hd__a21o_1
X_5380_ VPWR VGND VPWR VGND _1348_ _2108_ _1026_ _2112_ sky130_fd_sc_hd__or3_1
XFILLER_0_1_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4331_ VGND VPWR _1178_ _0656_ _1029_ i_tinyqv.cpu.alu_op\[0\] VPWR VGND sky130_fd_sc_hd__and3_1
X_4262_ VGND VPWR VPWR VGND _1109_ _1107_ _1108_ _1104_ sky130_fd_sc_hd__mux2_1
X_7050_ VPWR VGND VGND VPWR _2140_ _3329_ _3363_ sky130_fd_sc_hd__nor2_1
X_6001_ VGND VPWR _0267_ _2566_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4193_ VGND VPWR _1039_ _1040_ i_tinyqv.cpu.i_core.i_shift.b\[3\] VPWR VGND sky130_fd_sc_hd__xnor2_1
X_7952_ i_tinyqv.cpu.i_core.mcause\[4\] clknet_leaf_23_clk _0090_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_6903_ VGND VPWR _0476_ _3259_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7883_ i_tinyqv.cpu.i_core.i_registers.reg_access\[2\]\[2\] clknet_leaf_5_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[6\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6834_ VGND VPWR VPWR VGND _3206_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[28\]
+ net31 _0902_ sky130_fd_sc_hd__mux2_1
X_6765_ VPWR VGND VGND VPWR _3144_ _3029_ _3143_ sky130_fd_sc_hd__or2_1
X_3977_ VPWR VGND VGND VPWR _0708_ net79 _0829_ sky130_fd_sc_hd__nor2_1
X_5716_ VGND VPWR _0184_ _2365_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.i_regbuf\[28\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[28\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_8504_ i_tinyqv.cpu.i_core.i_instrret.register\[10\] clknet_leaf_49_clk i_tinyqv.cpu.i_core.i_instrret.reg_buf\[10\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_443 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6696_ VPWR VGND VGND VPWR _2991_ _3081_ _3080_ sky130_fd_sc_hd__nand2_1
X_8435_ i_tinyqv.cpu.imm\[13\] clknet_leaf_8_clk _0533_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_33_627 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5647_ VPWR VGND _2316_ i_tinyqv.cpu.instr_data_in\[8\] VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_0_5_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_5578_ VGND VPWR VGND VPWR _0144_ net241 _2263_ _2267_ _2240_ sky130_fd_sc_hd__o211a_1
X_8366_ i_tinyqv.cpu.instr_fetch_running clknet_leaf_22_clk _0465_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_4529_ VGND VPWR VGND VPWR _1368_ _0986_ _1366_ net4 _1367_ sky130_fd_sc_hd__a211o_1
Xhold241 net270 i_uart_tx.fsm_state\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_8297_ i_tinyqv.mem.q_ctrl.nibbles_remaining\[0\] clknet_leaf_14_clk _0396_ VPWR
+ VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold252 net281 i_tinyqv.cpu.instr_data\[3\]\[15\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold230 net259 i_tinyqv.cpu.imm\[12\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7317_ VPWR VGND VPWR VGND _3290_ _3374_ _3587_ _3556_ _3586_ _2149_ sky130_fd_sc_hd__a221o_1
Xhold274 net303 i_tinyqv.mem.q_ctrl.addr\[11\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 net314 i_tinyqv.cpu.data_addr\[11\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 net292 i_tinyqv.mem.data_from_read\[20\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7248_ VPWR VGND VGND VPWR net135 _3360_ _3529_ _0551_ sky130_fd_sc_hd__o21a_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.i_regbuf\[17\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[17\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[21\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7179_ VPWR VGND VGND VPWR _3478_ _3474_ net257 _3475_ _0533_ sky130_fd_sc_hd__o22a_1
XFILLER_0_36_421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_17_690 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_23_159 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xinput9 VGND VPWR net9 ui_in[7] VPWR VGND sky130_fd_sc_hd__buf_1
X_4880_ VGND VPWR VPWR VGND _1683_ i_tinyqv.cpu.debug_rd\[2\] _1680_ net150 sky130_fd_sc_hd__mux2_1
X_3900_ VPWR VGND _0752_ _0611_ VPWR VGND sky130_fd_sc_hd__buf_4
X_3831_ VPWR VGND VGND VPWR _0662_ _0661_ _0683_ _0660_ _0663_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_67_590 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6550_ VGND VPWR _0423_ _2959_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_3762_ VPWR VGND _0614_ i_tinyqv.cpu.counter\[3\] VPWR VGND sky130_fd_sc_hd__buf_4
XFILLER_0_6_304 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5501_ VGND VPWR _2209_ _2200_ _2213_ net214 VPWR VGND sky130_fd_sc_hd__o21ai_1
X_6481_ VGND VPWR _0413_ _2900_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_498 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_8220_ i_tinyqv.cpu.i_core.multiplier.accum\[3\] clknet_leaf_42_clk _0021_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5432_ VPWR VGND VPWR VGND _2159_ _1679_ _2147_ _2160_ sky130_fd_sc_hd__a21o_1
X_8151_ i_tinyqv.cpu.data_addr\[26\] clknet_leaf_35_clk _0263_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_5363_ VGND VPWR _1395_ _2097_ _2098_ _0788_ VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_321 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_4314_ VPWR VGND VPWR VGND _1156_ _1080_ _1160_ _1161_ sky130_fd_sc_hd__a21oi_1
X_7102_ VGND VPWR VPWR VGND _3411_ _3308_ _2126_ _3305_ _2132_ _1483_ sky130_fd_sc_hd__a32o_1
X_8082_ gpio_out_sel\[1\] clknet_leaf_19_clk _0009_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5294_ VGND VPWR VPWR VGND _2043_ _0018_ _2045_ sky130_fd_sc_hd__xor2_1
X_4245_ VPWR VGND _1092_ _1091_ VPWR VGND sky130_fd_sc_hd__buf_2
X_7033_ VPWR VGND VGND VPWR _1478_ _3337_ _3347_ sky130_fd_sc_hd__nor2_1
X_4176_ VPWR VGND VPWR VGND _1022_ i_tinyqv.cpu.i_core.load_top_bit _0878_ _1023_
+ sky130_fd_sc_hd__a21o_1
X_7935_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[26\] clknet_leaf_36_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[26\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_7866_ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[21\] clknet_leaf_53_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[21\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6817_ VPWR VGND VGND VPWR _1390_ _3191_ _2540_ sky130_fd_sc_hd__nand2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.i_regbuf\[29\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[29\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[1\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7797_ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[16\] clknet_leaf_3_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[16\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6748_ VGND VPWR VGND VPWR _3126_ _3128_ _3127_ sky130_fd_sc_hd__or2b_1
X_6679_ VPWR VGND VGND VPWR _3063_ _3065_ _3064_ sky130_fd_sc_hd__nand2_1
X_8418_ i_tinyqv.cpu.is_branch clknet_leaf_6_clk _0516_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_8349_ i_tinyqv.cpu.instr_data_start\[7\] clknet_leaf_36_clk _0448_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.i_regbuf\[18\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[18\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[22\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_53_clk VGND VPWR clknet_3_1__leaf_clk clknet_leaf_53_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.i_regbuf\[21\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[21\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[25\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.i_regbuf\[17\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[17\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[21\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_instrret.i_regbuf\[31\] i_tinyqv.cpu.i_core.i_instrret.reg_buf\[31\]
+ i_tinyqv.cpu.i_core.i_instrret.register\[3\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_cycles.i_regbuf\[15\] i_tinyqv.cpu.i_core.i_cycles.reg_buf\[15\]
+ i_tinyqv.cpu.i_core.i_cycles.register\[19\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_10_Right_10 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4030_ VPWR VGND _0852_ _0877_ _0849_ VPWR VGND sky130_fd_sc_hd__and2_2
X_5981_ VPWR VGND VPWR VGND _2552_ i_tinyqv.cpu.data_addr\[24\] _1758_ _2553_ i_tinyqv.cpu.i_core.i_shift.a\[28\]
+ sky130_fd_sc_hd__a22o_1
X_4932_ VGND VPWR VPWR VGND _1709_ uio_out[1] i_tinyqv.mem.q_ctrl.addr\[20\] _1716_
+ _1711_ _1712_ sky130_fd_sc_hd__a221o_4
X_7720_ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[3\] clknet_leaf_57_clk _0033_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_44_clk VGND VPWR clknet_3_5__leaf_clk clknet_leaf_44_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_7651_ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[30\] clknet_leaf_47_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[30\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6602_ VPWR VGND VPWR VGND i_tinyqv.cpu.i_core.imm_lo\[1\] _0749_ _2997_ _2999_ sky130_fd_sc_hd__a21oi_1
X_4863_ VGND VPWR VPWR VGND _1673_ i_tinyqv.cpu.debug_rd\[3\] _1669_ i_tinyqv.cpu.i_core.i_registers.reg_access\[9\]\[3\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA_14 i_tinyqv.cpu.i_core.mepc\[2\] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_4794_ VGND VPWR VGND VPWR _1629_ _0997_ _1628_ i_uart_rx.recieved_data\[3\] _0971_
+ sky130_fd_sc_hd__a211o_1
XANTENNA_47 i_tinyqv.cpu.i_core.imm_lo\[9\] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_0_6_112 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7582_ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[25\] clknet_leaf_58_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[25\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_3814_ _0666_ _0660_ _0661_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
XANTENNA_25 net69 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_36 i_tinyqv.cpu.i_core.imm_lo\[4\] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_6533_ VGND VPWR VPWR VGND _2944_ i_tinyqv.cpu.data_out\[19\] _2912_ i_tinyqv.cpu.data_out\[27\]
+ sky130_fd_sc_hd__mux2_1
X_6464_ VGND VPWR _2888_ _2832_ _2889_ net145 VPWR VGND sky130_fd_sc_hd__o21ai_1
X_5415_ VPWR VGND VPWR VGND _1510_ _2137_ _2145_ _2141_ _1460_ _2144_ sky130_fd_sc_hd__a221o_1
X_8203_ i_tinyqv.cpu.i_core.i_shift.a\[22\] clknet_leaf_40_clk _0315_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_6395_ VPWR VGND VPWR VGND _2833_ _2795_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5346_ VGND VPWR VPWR VGND _2085_ i_tinyqv.cpu.i_core.interrupt_req\[0\] _2084_ net250
+ sky130_fd_sc_hd__mux2_1
X_8134_ i_tinyqv.cpu.data_addr\[9\] clknet_leaf_32_clk _0246_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_8065_ i_spi.spi_clk_out clknet_leaf_27_clk _0200_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5277_ VPWR VGND VGND VPWR _2029_ _1975_ _2023_ sky130_fd_sc_hd__or2_1
X_4228_ VGND VPWR VPWR VGND _1075_ _1074_ _1058_ _1067_ sky130_fd_sc_hd__mux2_1
X_7016_ VPWR VGND VGND VPWR _2140_ _3295_ _3333_ sky130_fd_sc_hd__nor2_1
X_4159_ VGND VPWR VGND VPWR _1006_ _0997_ _1002_ i_uart_rx.recieved_data\[0\] _1005_
+ sky130_fd_sc_hd__a211o_1
Xmax_cap27 VGND VPWR net27 _0634_ VPWR VGND sky130_fd_sc_hd__buf_1
X_7918_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[9\] clknet_leaf_24_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[9\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_35_clk VGND VPWR clknet_3_7__leaf_clk clknet_leaf_35_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_7849_ i_tinyqv.cpu.i_core.i_registers.reg_access\[5\]\[0\] clknet_leaf_45_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[4\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_273 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_21_449 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.i_regbuf\[22\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[22\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[26\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.i_regbuf\[29\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[29\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[1\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_26_clk VGND VPWR clknet_3_6__leaf_clk clknet_leaf_26_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_0_29_505 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xinput12 VGND VPWR net12 uio_in[4] VPWR VGND sky130_fd_sc_hd__buf_1
X_5200_ VPWR VGND VGND VPWR _1955_ _1902_ _1950_ sky130_fd_sc_hd__or2_1
X_6180_ VGND VPWR VPWR VGND _2671_ i_tinyqv.cpu.i_core.mepc\[17\] _2667_ i_tinyqv.cpu.i_core.mepc\[13\]
+ sky130_fd_sc_hd__mux2_1
X_5131_ VPWR VGND VGND VPWR _1887_ _1889_ _1888_ sky130_fd_sc_hd__nand2_1
X_5062_ _1823_ _1797_ _1799_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_4013_ VPWR VGND VGND VPWR net127 _0837_ _0863_ _0029_ sky130_fd_sc_hd__o21a_1
XFILLER_0_75_600 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_17_clk VGND VPWR clknet_3_3__leaf_clk clknet_leaf_17_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_5964_ VGND VPWR _0255_ _2541_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7703_ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[18\] clknet_leaf_53_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[18\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5895_ VGND VPWR VPWR VGND _2494_ i_spi.data\[4\] _2386_ i_debug_uart_tx.uart_tx_data\[5\]
+ sky130_fd_sc_hd__mux2_1
X_4915_ VGND VPWR VPWR VGND _1703_ _1303_ _1701_ net268 sky130_fd_sc_hd__mux2_1
X_4846_ VGND VPWR _0037_ _1663_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7634_ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[13\] clknet_leaf_55_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[13\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7565_ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[8\] clknet_leaf_57_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[8\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.i_regbuf\[10\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[10\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[14\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6516_ VGND VPWR VGND VPWR _2929_ _2906_ _0864_ sky130_fd_sc_hd__xnor2_4
X_4777_ VPWR VGND VPWR VGND _1606_ _1612_ _1611_ i_tinyqv.cpu.i_core.i_instrret.data\[3\]
+ _0929_ _1608_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_70_360 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7496_ VPWR VGND VGND VPWR _3733_ _3234_ _3239_ _3732_ _3734_ sky130_fd_sc_hd__o22a_1
XFILLER_0_43_574 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6447_ VGND VPWR _0403_ _2876_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_660 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_6378_ VGND VPWR VPWR VGND _2818_ _2817_ _2800_ _2816_ sky130_fd_sc_hd__mux2_1
X_8117_ i_tinyqv.cpu.instr_data\[3\]\[1\] clknet_leaf_9_clk _0229_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_482 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_5329_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_cycles.cy _0744_ i_tinyqv.cpu.i_core.cycle_count\[0\]
+ _2071_ sky130_fd_sc_hd__o21a_1
X_8048_ i_debug_uart_tx.cycle_counter\[2\] clknet_leaf_30_clk _0183_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.i_regbuf\[7\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[7\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[11\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_129 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_28_25 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_44_79 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5680_ VPWR VGND _2341_ _2340_ VPWR VGND sky130_fd_sc_hd__buf_2
X_4700_ VGND VPWR VGND VPWR _1536_ i_tinyqv.cpu.data_read_n\[1\] i_tinyqv.cpu.data_read_n\[0\]
+ i_tinyqv.cpu.data_write_n\[1\] i_tinyqv.cpu.data_write_n\[0\] _0865_ sky130_fd_sc_hd__a41o_2
XFILLER_0_17_519 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.i_regbuf\[5\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[5\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[9\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4631_ VPWR VGND VGND VPWR _1448_ _1467_ _1466_ sky130_fd_sc_hd__nand2_1
X_4562_ VGND VPWR VGND VPWR _1387_ _1398_ _1397_ sky130_fd_sc_hd__and2_4
X_7350_ VPWR VGND VPWR VGND _3611_ _3612_ _1439_ _3613_ sky130_fd_sc_hd__or3_1
X_6301_ VGND VPWR VPWR VGND _2760_ _1721_ _1552_ net256 sky130_fd_sc_hd__mux2_1
X_4493_ VPWR VGND VPWR VGND _1280_ _1030_ _1331_ _1332_ sky130_fd_sc_hd__a21o_1
X_7281_ VPWR VGND _3558_ _3554_ _3299_ _3291_ _3557_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_6232_ VPWR VGND VGND VPWR _2041_ _2712_ _2711_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_6_clk VGND VPWR clknet_3_1__leaf_clk clknet_leaf_6_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_0_0_641 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_6163_ VGND VPWR VPWR VGND _2662_ i_tinyqv.cpu.i_core.mepc\[9\] _2656_ i_tinyqv.cpu.i_core.mepc\[5\]
+ sky130_fd_sc_hd__mux2_1
X_5114_ VPWR VGND _1873_ _1872_ _1871_ VPWR VGND sky130_fd_sc_hd__and2_1
X_6094_ VGND VPWR VPWR VGND _2615_ i_tinyqv.cpu.i_core.i_shift.a\[19\] _2595_ i_tinyqv.cpu.i_core.i_shift.a\[23\]
+ sky130_fd_sc_hd__mux2_1
X_5045_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[3\] _1806_ _1789_ sky130_fd_sc_hd__nand2_1
X_6996_ VPWR VGND VPWR VGND _3317_ _3304_ _3312_ _3315_ _3316_ _3282_ sky130_fd_sc_hd__o32a_1
X_5947_ VGND VPWR VPWR VGND _2530_ i_tinyqv.cpu.i_core.mepc\[13\] _2106_ i_tinyqv.cpu.i_core.i_shift.a\[17\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_485 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5878_ VGND VPWR _0227_ _2483_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7617_ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[28\] clknet_leaf_0_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[28\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.i_regbuf\[11\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[11\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[15\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4829_ VGND VPWR VPWR VGND _1654_ i_tinyqv.cpu.debug_rd\[0\] _1653_ net215 sky130_fd_sc_hd__mux2_1
X_7548_ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[23\] clknet_leaf_46_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[23\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7479_ VPWR VGND VGND VPWR _3719_ i_tinyqv.cpu.instr_data_start\[21\] _3715_ sky130_fd_sc_hd__or2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.i_regbuf\[4\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[4\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[8\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_34_393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6850_ VPWR VGND VPWR VGND i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[29\] _2987_
+ _3221_ _2306_ _1211_ _3028_ sky130_fd_sc_hd__a221o_1
X_5801_ VGND VPWR VGND VPWR _0204_ net97 _2427_ _2430_ _2221_ sky130_fd_sc_hd__o211a_1
X_6781_ VGND VPWR _3157_ _3158_ _3155_ VPWR VGND sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_8_Right_8 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5732_ VGND VPWR _0188_ _2377_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8520_ i_tinyqv.cpu.i_core.i_instrret.register\[26\] clknet_leaf_50_clk i_tinyqv.cpu.i_core.i_instrret.reg_buf\[26\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_3993_ VPWR VGND VPWR VGND _0844_ i_tinyqv.cpu.alu_op\[1\] sky130_fd_sc_hd__inv_2
X_5663_ VGND VPWR VPWR VGND _2326_ _1720_ _2308_ i_tinyqv.cpu.instr_data\[3\]\[14\]
+ sky130_fd_sc_hd__mux2_1
X_8451_ i_tinyqv.cpu.imm\[29\] clknet_leaf_22_clk _0549_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5594_ VPWR VGND VGND VPWR _2278_ i_uart_rx.rxd_reg\[0\] _2276_ sky130_fd_sc_hd__or2_1
X_8382_ i_debug_uart_tx.uart_tx_data\[7\] clknet_leaf_19_clk _0480_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
X_7402_ VGND VPWR VPWR VGND _3655_ net312 _3624_ i_tinyqv.mem.q_ctrl.addr\[4\] sky130_fd_sc_hd__mux2_1
X_4614_ VGND VPWR VPWR VGND _1450_ i_tinyqv.cpu.instr_data\[3\]\[5\] _1449_ i_tinyqv.cpu.instr_data\[1\]\[5\]
+ sky130_fd_sc_hd__mux2_1
X_4545_ VGND VPWR VPWR VGND _1382_ debug_rd_r\[1\] debug_register_data i_spi.data\[7\]
+ sky130_fd_sc_hd__mux2_1
X_7333_ VGND VPWR _0565_ _3600_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4476_ VPWR VGND VPWR VGND _1310_ _1315_ _1311_ _1313_ sky130_fd_sc_hd__or3b_2
X_7264_ VGND VPWR _0553_ _3543_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_396 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6215_ VPWR VGND VGND VPWR _2695_ _1999_ _2694_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_39_Right_39 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7195_ VPWR VGND VPWR VGND _3491_ _3476_ _3479_ _3492_ sky130_fd_sc_hd__a21o_1
X_6146_ VGND VPWR VPWR VGND _2652_ _2651_ _2645_ i_tinyqv.cpu.i_core.i_shift.b\[2\]
+ sky130_fd_sc_hd__mux2_1
X_6077_ VGND VPWR _0303_ _2606_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5028_ VPWR VGND VPWR VGND i_tinyqv.cpu.i_core.i_shift.a\[2\] _1789_ _1790_ i_tinyqv.cpu.i_core.i_shift.a\[3\]
+ _1309_ sky130_fd_sc_hd__a22oi_1
X_6979_ VPWR VGND VGND VPWR _3299_ _3300_ _3301_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_48_Right_48 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_51_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_360 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_57_Right_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_66_Right_66 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.i_regbuf\[11\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[11\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[15\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_157 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_75_Right_75 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_10_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_4330_ VPWR VGND VGND VPWR _1030_ _1177_ _0919_ sky130_fd_sc_hd__nand2_1
X_4261_ VGND VPWR i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt\[1\] _1108_ VPWR
+ VGND sky130_fd_sc_hd__clkbuf_4
X_6000_ VGND VPWR VPWR VGND _2566_ i_tinyqv.cpu.instr_data\[2\]\[4\] _2563_ i_tinyqv.cpu.instr_data_in\[4\]
+ sky130_fd_sc_hd__mux2_1
X_4192_ VGND VPWR _1027_ _1039_ _0907_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_7951_ i_tinyqv.cpu.i_core.mcause\[3\] clknet_leaf_38_clk _0089_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_6902_ VGND VPWR VPWR VGND _3259_ _2631_ _3254_ i_debug_uart_tx.uart_tx_data\[3\]
+ sky130_fd_sc_hd__mux2_1
X_7882_ i_tinyqv.cpu.i_core.i_registers.reg_access\[2\]\[1\] clknet_leaf_5_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[5\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6833_ VGND VPWR VGND VPWR _0460_ i_tinyqv.cpu.instr_data_start\[19\] _3123_ _3204_
+ _3205_ sky130_fd_sc_hd__o211a_1
X_6764_ VGND VPWR VPWR VGND _3143_ _3142_ _3047_ _3135_ sky130_fd_sc_hd__mux2_1
X_3976_ VPWR VGND VGND VPWR _0799_ _0815_ _0828_ sky130_fd_sc_hd__nor2_1
X_5715_ VGND VPWR _2365_ _2363_ _2357_ _2364_ VPWR VGND sky130_fd_sc_hd__and3_1
X_6695_ VGND VPWR VPWR VGND _3078_ _3080_ _3079_ sky130_fd_sc_hd__xor2_1
X_8503_ i_tinyqv.cpu.i_core.i_instrret.register\[9\] clknet_leaf_45_clk i_tinyqv.cpu.i_core.i_instrret.reg_buf\[9\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_455 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_8434_ i_tinyqv.cpu.imm\[12\] clknet_leaf_8_clk _0532_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_5646_ VGND VPWR _0164_ _2315_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_488 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_60_436 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5577_ VPWR VGND VGND VPWR _2267_ i_uart_rx.recieved_data\[2\] _2264_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_149 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold220 net249 i_tinyqv.cpu.is_alu_imm VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_8365_ i_tinyqv.cpu.instr_data_start\[23\] clknet_leaf_36_clk _0464_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
Xhold242 net271 i_tinyqv.mem.q_ctrl.spi_in_buffer\[6\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4528_ VPWR VGND VPWR VGND _1001_ i_spi.data\[2\] _1000_ _1367_ uo_out[2] sky130_fd_sc_hd__a22o_1
Xhold253 net282 i_spi.spi_dc VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_8296_ i_tinyqv.mem.q_ctrl.data_req clknet_leaf_16_clk _0395_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_2
Xhold231 net260 i_tinyqv.cpu.instr_data\[3\]\[3\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7316_ VPWR VGND VGND VPWR _3313_ _3586_ _3454_ sky130_fd_sc_hd__nand2_1
Xhold275 net304 i_tinyqv.mem.q_ctrl.addr\[13\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 net315 i_tinyqv.mem.q_ctrl.addr\[14\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 net293 i_tinyqv.mem.qspi_data_buf\[12\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4459_ VGND VPWR VGND VPWR _1302_ _1252_ _1261_ _0846_ _1301_ sky130_fd_sc_hd__a211o_1
X_7247_ VGND VPWR VGND VPWR _3529_ _3464_ _3499_ _3328_ _3438_ sky130_fd_sc_hd__a211o_1
X_7178_ VGND VPWR VPWR VGND _3478_ _3476_ _2123_ _3328_ _3331_ _2155_ sky130_fd_sc_hd__a32o_1
X_6129_ VPWR VGND VGND VPWR _2638_ _1400_ i_tinyqv.cpu.instr_data\[0\]\[1\] sky130_fd_sc_hd__or2_1
XFILLER_0_68_558 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_36_14 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_36_25 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_3830_ VPWR VGND VPWR VGND _0681_ i_tinyqv.cpu.i_core.i_registers.reg_access\[9\]\[3\]
+ _0680_ _0682_ i_tinyqv.cpu.i_core.i_registers.reg_access\[6\]\[3\] sky130_fd_sc_hd__a22o_1
X_3761_ VPWR VGND VGND VPWR _0612_ _0613_ _0611_ sky130_fd_sc_hd__nor2_2
X_5500_ VPWR VGND _2212_ _2209_ i_uart_tx.cycle_counter\[6\] VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_54_241 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_6480_ VGND VPWR VPWR VGND _2900_ i_tinyqv.mem.q_ctrl.spi_in_buffer\[2\] _2897_ net12
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_5431_ VPWR VGND VPWR VGND i_tinyqv.cpu.i_core.i_registers.rd\[0\] i_tinyqv.cpu.i_core.i_registers.rd\[1\]
+ i_tinyqv.cpu.i_core.i_registers.rd\[2\] _2159_ sky130_fd_sc_hd__a21o_1
X_8150_ i_tinyqv.cpu.data_addr\[25\] clknet_leaf_40_clk _0262_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_5362_ VGND VPWR VGND VPWR _2097_ net18 _2096_ _0798_ _2056_ sky130_fd_sc_hd__a211o_1
X_8081_ gpio_out_sel\[0\] clknet_leaf_19_clk _0008_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4313_ VPWR VGND VPWR VGND _1159_ _1091_ _1076_ _1160_ sky130_fd_sc_hd__a21o_1
X_7101_ VPWR VGND VGND VPWR _3410_ _3287_ _3352_ _3337_ _3292_ _1478_ sky130_fd_sc_hd__o41a_1
X_5293_ VPWR VGND VGND VPWR _2017_ _2045_ _2044_ sky130_fd_sc_hd__nand2_1
X_7032_ VPWR VGND VGND VPWR _2120_ _2130_ _3346_ sky130_fd_sc_hd__nor2_1
X_4244_ VPWR VGND VGND VPWR _1091_ _1042_ _1057_ sky130_fd_sc_hd__nand2_2
X_4175_ VPWR VGND VPWR VGND _1022_ _0955_ sky130_fd_sc_hd__inv_2
X_7934_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[25\] clknet_leaf_24_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[25\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7865_ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[20\] clknet_leaf_48_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[20\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6816_ VGND VPWR _3189_ _3190_ _3186_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_7796_ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[15\] clknet_leaf_0_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[15\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6747_ VPWR VGND VGND VPWR _0726_ _3127_ i_tinyqv.cpu.imm\[12\] sky130_fd_sc_hd__nand2_1
X_3959_ VPWR VGND VPWR VGND _0619_ i_tinyqv.cpu.imm\[14\] _0617_ _0811_ i_tinyqv.cpu.i_core.imm_lo\[6\]
+ sky130_fd_sc_hd__a22o_1
X_6678_ VPWR VGND VGND VPWR _3064_ _0883_ i_tinyqv.cpu.i_core.imm_lo\[6\] sky130_fd_sc_hd__or2_1
X_5629_ VPWR VGND VPWR VGND _2305_ _2304_ sky130_fd_sc_hd__inv_2
X_8417_ i_tinyqv.cpu.is_lui clknet_leaf_7_clk _0515_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_8348_ i_tinyqv.cpu.instr_data_start\[6\] clknet_leaf_24_clk _0447_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_8279_ i_tinyqv.mem.data_from_read\[19\] clknet_leaf_21_clk _0378_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.i_regbuf\[25\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[25\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[29\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_377 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.i_regbuf\[14\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[14\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[18\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_instrret.i_regbuf\[24\] i_tinyqv.cpu.i_core.i_instrret.reg_buf\[24\]
+ i_tinyqv.cpu.i_core.i_instrret.register\[28\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_2_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_5980_ VPWR VGND VGND VPWR _2107_ _1758_ _2552_ sky130_fd_sc_hd__nor2_1
X_4931_ VPWR VGND VGND VPWR _1715_ i_tinyqv.mem.q_ctrl.nibbles_remaining\[0\] _1713_
+ _1716_ sky130_fd_sc_hd__nor3_1
XFILLER_0_59_355 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_4862_ VGND VPWR _0080_ _1672_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7650_ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[29\] clknet_leaf_58_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[29\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6601_ VGND VPWR _2998_ i_tinyqv.cpu.i_core.imm_lo\[1\] _0749_ _2997_ VPWR VGND sky130_fd_sc_hd__and3_1
X_3813_ VGND VPWR VGND VPWR _0664_ _0630_ _0659_ _0665_ i_tinyqv.cpu.i_core.i_registers.reg_access\[11\]\[3\]
+ sky130_fd_sc_hd__a2bb2o_1
X_4793_ VPWR VGND VPWR VGND i_spi.data\[3\] _1000_ _1628_ _0986_ net5 _1627_ sky130_fd_sc_hd__a221o_1
XFILLER_0_55_561 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XANTENNA_15 i_tinyqv.cpu.imm\[14\] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_7581_ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[24\] clknet_leaf_59_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[24\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XANTENNA_26 _1302_ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_37 i_tinyqv.cpu.i_core.imm_lo\[9\] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_48 i_tinyqv.cpu.i_core.imm_lo\[9\] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_6532_ VGND VPWR _0421_ _2943_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_669 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_15_425 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6463_ VGND VPWR VGND VPWR _2888_ _2797_ _2803_ _2842_ _2887_ sky130_fd_sc_hd__o211a_1
X_8202_ i_tinyqv.cpu.i_core.i_shift.a\[21\] clknet_leaf_40_clk _0314_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5414_ VPWR VGND VPWR VGND _1478_ _2118_ _2144_ _2135_ _2142_ _2143_ sky130_fd_sc_hd__a221o_1
X_6394_ VPWR VGND _2832_ _2304_ VPWR VGND sky130_fd_sc_hd__buf_2
X_8133_ i_tinyqv.cpu.data_addr\[8\] clknet_leaf_32_clk _0245_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_5345_ VPWR VGND VGND VPWR _2081_ _2083_ _2084_ sky130_fd_sc_hd__nor2_1
X_8064_ i_spi.spi_select clknet_leaf_26_clk net185 VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5276_ VPWR VGND _2028_ _2027_ _2026_ VPWR VGND sky130_fd_sc_hd__and2_1
X_4227_ VGND VPWR VPWR VGND _1074_ _1073_ i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt\[1\]
+ _1070_ sky130_fd_sc_hd__mux2_1
X_7015_ VGND VPWR VGND VPWR _0515_ net212 _3282_ _3332_ _1753_ sky130_fd_sc_hd__o211a_1
X_4158_ VPWR VGND VPWR VGND _1004_ gpio_out_sel\[0\] _1003_ _1005_ i_spi.busy sky130_fd_sc_hd__a22o_1
XFILLER_0_69_108 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4089_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.imm_lo\[4\] i_tinyqv.cpu.i_core.imm_lo\[5\]
+ i_tinyqv.cpu.i_core.imm_lo\[7\] _0936_ sky130_fd_sc_hd__nor3_1
X_7917_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[8\] clknet_leaf_39_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[8\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7848_ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[3\] clknet_leaf_50_clk _0069_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7779_ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[30\] clknet_leaf_54_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[30\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.i_regbuf\[30\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[30\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[2\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_200 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.i_regbuf\[26\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[26\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[30\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.i_regbuf\[15\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[15\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[19\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_517 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xinput13 VGND VPWR net13 uio_in[5] VPWR VGND sky130_fd_sc_hd__buf_1
X_5130_ VPWR VGND VGND VPWR _1888_ i_tinyqv.cpu.i_core.multiplier.accum\[9\] _1886_
+ sky130_fd_sc_hd__or2_1
X_5061_ VGND VPWR VPWR VGND _1820_ _1822_ _1821_ sky130_fd_sc_hd__xor2_1
X_4012_ VPWR VGND VPWR VGND _0863_ _0862_ sky130_fd_sc_hd__inv_2
X_5963_ VGND VPWR VPWR VGND _2541_ _2540_ _2524_ i_tinyqv.cpu.data_addr\[18\] sky130_fd_sc_hd__mux2_1
X_7702_ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[17\] clknet_leaf_56_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[17\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4914_ VGND VPWR _0054_ _1702_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5894_ VGND VPWR _0233_ _2493_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_325 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7633_ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[12\] clknet_leaf_56_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[12\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4845_ VGND VPWR VPWR VGND _1663_ i_tinyqv.cpu.debug_rd\[3\] _1659_ i_tinyqv.cpu.i_core.i_registers.reg_access\[11\]\[3\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_317 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7564_ i_tinyqv.cpu.i_core.i_registers.reg_access\[14\]\[3\] clknet_leaf_57_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[7\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4776_ VPWR VGND VPWR VGND net15 _0991_ _1611_ _1609_ i_tinyqv.cpu.i_core.mstatus_mpie
+ _1610_ sky130_fd_sc_hd__a221o_1
X_6515_ VGND VPWR VPWR VGND _2928_ i_spi.dc_in _2909_ i_debug_uart_tx.uart_tx_data\[1\]
+ sky130_fd_sc_hd__mux2_1
X_7495_ VPWR VGND VPWR VGND _3726_ i_tinyqv.cpu.instr_data_start\[23\] i_tinyqv.cpu.was_early_branch
+ _3733_ sky130_fd_sc_hd__a21o_1
X_6446_ _2876_ _2806_ _2792_ _2811_ _2875_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.i_regbuf\[8\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[8\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[12\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6377_ VGND VPWR VPWR VGND _2817_ _2815_ _2797_ i_tinyqv.mem.q_ctrl.delay_cycles_cfg\[1\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_160 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_8116_ i_tinyqv.cpu.instr_data\[3\]\[0\] clknet_leaf_9_clk _0228_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5328_ VPWR VGND VPWR VGND _1026_ net99 _2070_ _0091_ sky130_fd_sc_hd__a21o_1
X_8047_ i_debug_uart_tx.cycle_counter\[1\] clknet_leaf_30_clk _0182_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5259_ VPWR VGND VGND VPWR _1981_ _1984_ _2012_ _2010_ sky130_fd_sc_hd__nand3_1
XFILLER_0_26_509 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_34_542 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_61_372 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_1_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.i_regbuf\[7\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[7\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[11\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_24 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_56_177 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4630_ _1456_ _1460_ _1466_ _1465_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_6300_ VGND VPWR _0373_ _2759_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4561_ VGND VPWR _1396_ _1389_ _1397_ _1391_ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_4492_ VGND VPWR _1299_ _1125_ _1331_ _1030_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_7280_ VGND VPWR VPWR VGND _3557_ _3556_ _3555_ _2165_ _3337_ _2123_ sky130_fd_sc_hd__a32o_1
X_6231_ VGND VPWR VGND VPWR _2711_ _2044_ _2017_ _2043_ sky130_fd_sc_hd__a21bo_1
X_6162_ VGND VPWR _0333_ _2661_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5113_ VPWR VGND VGND VPWR _1872_ _1868_ _1870_ sky130_fd_sc_hd__or2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.i_regbuf\[5\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[5\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[9\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_697 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6093_ VGND VPWR _0311_ _2614_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5044_ VGND VPWR _1805_ _0019_ _1787_ VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_6995_ VPWR VGND VPWR VGND _3316_ i_tinyqv.cpu.is_auipc sky130_fd_sc_hd__inv_2
X_5946_ VGND VPWR _0249_ _2529_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5877_ VGND VPWR VPWR VGND _2483_ net283 _2468_ _1721_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_689 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_7616_ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[27\] clknet_leaf_2_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[27\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4828_ VGND VPWR VGND VPWR _1653_ _1189_ _1640_ i_tinyqv.cpu.i_core.i_registers.rd\[1\]
+ sky130_fd_sc_hd__and3b_2
XFILLER_0_47_177 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4759_ VGND VPWR VGND VPWR _0748_ _0612_ _1591_ _1594_ _1593_ sky130_fd_sc_hd__a2bb2o_1
X_7547_ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[22\] clknet_leaf_46_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[22\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_575 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_512 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_7478_ VPWR VGND VPWR VGND _3717_ _2733_ _3713_ _0592_ _3718_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_534 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_6429_ VGND VPWR _2861_ _2855_ _2862_ _2810_ VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_556 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.i_regbuf\[4\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[4\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[8\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_689 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5800_ VPWR VGND VPWR VGND _1725_ _1004_ net204 _2430_ sky130_fd_sc_hd__a21o_1
X_6780_ VPWR VGND VGND VPWR _3147_ _3156_ _3157_ sky130_fd_sc_hd__nor2_1
X_3992_ VPWR VGND VPWR VGND _0843_ i_tinyqv.cpu.alu_op\[2\] sky130_fd_sc_hd__inv_2
X_5731_ _2375_ _2376_ _2377_ _1729_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_5662_ VGND VPWR _0170_ _2325_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8450_ i_tinyqv.cpu.imm\[28\] clknet_leaf_9_clk _0548_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5593_ VPWR VGND VPWR VGND _2277_ _2276_ sky130_fd_sc_hd__inv_2
X_8381_ i_debug_uart_tx.uart_tx_data\[6\] clknet_leaf_19_clk _0479_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_7401_ VPWR VGND VGND VPWR i_tinyqv.cpu.data_addr\[8\] _2682_ _3005_ _3654_ sky130_fd_sc_hd__o21a_1
X_4613_ VGND VPWR _1414_ _1449_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_4544_ VGND VPWR _0052_ _1381_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7332_ VGND VPWR VPWR VGND _3600_ _0660_ _2153_ _3599_ sky130_fd_sc_hd__mux2_1
X_7263_ VGND VPWR VPWR VGND _3543_ _3542_ _3395_ _0656_ sky130_fd_sc_hd__mux2_1
X_4475_ VPWR VGND VGND VPWR _1311_ _1313_ _1314_ sky130_fd_sc_hd__nor2_1
X_6214_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[13\] _2694_ _1813_ sky130_fd_sc_hd__nand2_1
X_7194_ VPWR VGND VPWR VGND i_tinyqv.cpu.instr_data\[0\]\[0\] _3487_ _3491_ _3488_
+ i_tinyqv.cpu.instr_data\[1\]\[0\] _3490_ sky130_fd_sc_hd__a221o_1
X_6145_ VPWR VGND VPWR VGND _2651_ _2650_ sky130_fd_sc_hd__inv_2
X_6076_ VGND VPWR VPWR VGND _2606_ i_tinyqv.cpu.i_core.i_shift.a\[14\] _2593_ i_tinyqv.cpu.i_core.i_shift.a\[10\]
+ sky130_fd_sc_hd__mux2_1
X_5027_ VGND VPWR VPWR VGND _1789_ _0636_ _0641_ net73 i_tinyqv.cpu.i_core.cycle\[0\]
+ sky130_fd_sc_hd__o31a_2
X_6978_ VPWR VGND VGND VPWR _1498_ _3300_ _3287_ sky130_fd_sc_hd__nand2_1
X_5929_ VGND VPWR VPWR VGND _2518_ _2517_ _2502_ i_tinyqv.cpu.data_addr\[7\] sky130_fd_sc_hd__mux2_1
XFILLER_0_0_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_48_464 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_63_445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xsplit40 VPWR VGND net69 i_tinyqv.cpu.alu_op\[0\] VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_0_66_283 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4260_ VGND VPWR VPWR VGND _1107_ _1106_ _1103_ _1105_ sky130_fd_sc_hd__mux2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.i_regbuf\[29\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[29\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[1\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4191_ VPWR VGND VGND VPWR _1038_ i_tinyqv.cpu.i_core.i_shift.b\[4\] _1037_ sky130_fd_sc_hd__or2_1
X_7950_ i_tinyqv.cpu.i_core.mcause\[1\] clknet_leaf_38_clk _0088_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_6901_ VGND VPWR _0475_ _3258_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7881_ i_tinyqv.cpu.i_core.i_registers.reg_access\[2\]\[0\] clknet_leaf_49_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[4\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6832_ VGND VPWR _1752_ _3205_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_6763_ VGND VPWR VPWR VGND _3142_ _3141_ _2990_ _2530_ sky130_fd_sc_hd__mux2_1
X_3975_ VPWR VGND _0827_ _0815_ _0799_ VPWR VGND sky130_fd_sc_hd__and2_1
X_5714_ VPWR VGND VGND VPWR i_debug_uart_tx.cycle_counter\[3\] _2364_ _2360_ sky130_fd_sc_hd__nand2_1
X_6694_ VGND VPWR _3066_ _3063_ _3079_ _3065_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_8502_ i_tinyqv.cpu.i_core.i_instrret.register\[8\] clknet_leaf_49_clk i_tinyqv.cpu.i_core.i_instrret.reg_buf\[8\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_17_Left_98 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5645_ VGND VPWR VPWR VGND _2315_ i_tinyqv.cpu.instr_data_in\[7\] _2309_ i_tinyqv.cpu.instr_data\[3\]\[7\]
+ sky130_fd_sc_hd__mux2_1
X_8433_ i_tinyqv.cpu.i_core.imm_lo\[11\] clknet_leaf_22_clk _0531_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
X_5576_ VGND VPWR VGND VPWR _0143_ net225 _2263_ _2266_ _2240_ sky130_fd_sc_hd__o211a_1
Xhold210 net239 i_spi.bits_remaining\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_353 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_8364_ i_tinyqv.cpu.instr_data_start\[22\] clknet_leaf_36_clk _0463_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
X_8295_ i_tinyqv.mem.q_ctrl.read_cycles_count\[2\] clknet_leaf_15_clk _0394_ VPWR
+ VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4527_ VPWR VGND VPWR VGND i_uart_rx.recieved_data\[2\] _0996_ _1366_ net14 gpio_out_sel\[2\]
+ _0974_ sky130_fd_sc_hd__a221o_1
Xhold232 net261 i_tinyqv.mem.qspi_data_buf\[31\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 net250 i_tinyqv.cpu.i_core.last_interrupt_req\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 net272 i_tinyqv.cpu.instr_data\[3\]\[13\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7315_ VGND VPWR VPWR VGND _0662_ _3585_ i_tinyqv.cpu.mem_op_increment_reg sky130_fd_sc_hd__xor2_1
Xhold287 net316 i_debug_uart_tx.uart_tx_data\[6\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 net305 i_tinyqv.mem.q_ctrl.addr\[5\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 net294 i_tinyqv.cpu.data_write_n\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 net283 i_tinyqv.cpu.instr_data\[0\]\[15\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4458_ VGND VPWR VGND VPWR _1301_ _1030_ _1280_ _1300_ _1125_ sky130_fd_sc_hd__o211a_1
X_7246_ VGND VPWR _0550_ _3528_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7177_ VPWR VGND VGND VPWR _3477_ _3474_ net259 _3475_ _0532_ sky130_fd_sc_hd__o22a_1
X_4389_ VPWR VGND VPWR VGND i_spi.data\[5\] _1000_ _1232_ _0997_ i_uart_rx.recieved_data\[5\]
+ _0908_ sky130_fd_sc_hd__a221o_1
X_6128_ VGND VPWR _0323_ _2637_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6059_ VGND VPWR _0294_ _2597_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_3760_ VGND VPWR VGND VPWR _0608_ i_tinyqv.cpu.counter\[3\] _0612_ sky130_fd_sc_hd__or2_4
XFILLER_0_42_404 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5430_ VGND VPWR _0105_ _2158_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_2_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_5361_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.mepc\[2\] net18 _2096_ sky130_fd_sc_hd__nor2_1
X_8080_ i_uart_tx.txd_reg clknet_leaf_29_clk _0211_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5292_ VGND VPWR VGND VPWR _2044_ _2020_ _1993_ _2019_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_2_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_4312_ VGND VPWR VPWR VGND _1159_ _1158_ i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt\[1\]
+ _1157_ sky130_fd_sc_hd__mux2_1
X_7100_ VGND VPWR VPWR VGND _3409_ _3408_ _3319_ _3287_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_345 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4243_ VPWR VGND VGND VPWR _1080_ _1090_ _1089_ sky130_fd_sc_hd__nand2_1
X_7031_ VGND VPWR VGND VPWR _0518_ i_tinyqv.cpu.is_jal _3282_ _3345_ _1753_ sky130_fd_sc_hd__o211a_1
X_4174_ VPWR VGND VPWR VGND _0981_ _0956_ _1020_ _1021_ sky130_fd_sc_hd__a21o_1
X_7933_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[24\] clknet_leaf_37_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[24\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_345 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7864_ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[19\] clknet_leaf_48_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[19\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6815_ VGND VPWR VGND VPWR _3187_ _3189_ _3188_ sky130_fd_sc_hd__or2b_1
X_7795_ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[14\] clknet_leaf_56_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[14\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_710 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6746_ VPWR VGND VGND VPWR _0726_ i_tinyqv.cpu.imm\[12\] _3126_ sky130_fd_sc_hd__nor2_1
X_3958_ VPWR VGND VPWR VGND i_tinyqv.cpu.imm\[18\] _0615_ _0810_ _0617_ i_tinyqv.cpu.imm\[30\]
+ _0809_ sky130_fd_sc_hd__a221o_1
X_6677_ VPWR VGND VGND VPWR _0883_ _3063_ i_tinyqv.cpu.i_core.imm_lo\[6\] sky130_fd_sc_hd__nand2_1
X_3889_ VPWR VGND VGND VPWR net20 _0741_ _0740_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_426 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5628_ i_tinyqv.mem.q_ctrl.stop_txn_reg _2303_ _2304_ i_debug_uart_tx.resetn VGND
+ VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_8416_ i_tinyqv.cpu.is_alu_reg clknet_leaf_6_clk _0514_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5559_ VGND VPWR _2253_ _2242_ _2255_ i_uart_rx.cycle_counter\[7\] VPWR VGND sky130_fd_sc_hd__o21ai_1
X_8347_ i_tinyqv.cpu.instr_data_start\[5\] clknet_leaf_24_clk _0446_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.i_regbuf\[22\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[22\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[26\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_183 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_8278_ i_tinyqv.mem.data_from_read\[18\] clknet_leaf_17_clk _0377_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_7229_ VGND VPWR VPWR VGND _3518_ _3517_ _3396_ i_tinyqv.cpu.imm\[24\] sky130_fd_sc_hd__mux2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.i_regbuf\[18\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[18\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[22\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_instrret.i_regbuf\[17\] i_tinyqv.cpu.i_core.i_instrret.reg_buf\[17\]
+ i_tinyqv.cpu.i_core.i_instrret.register\[21\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4930_ VPWR VGND VGND VPWR _1715_ _1706_ _1714_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_304 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4861_ VGND VPWR VPWR VGND _1672_ i_tinyqv.cpu.debug_rd\[2\] _1669_ i_tinyqv.cpu.i_core.i_registers.reg_access\[9\]\[2\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_710 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6600_ VGND VPWR VPWR VGND net85 _2997_ i_tinyqv.cpu.i_core.imm_lo\[2\] sky130_fd_sc_hd__xor2_1
X_3812_ VGND VPWR _0662_ _0660_ _0664_ _0663_ _0661_ VPWR VGND sky130_fd_sc_hd__and4b_1
XPHY_EDGE_ROW_25_Left_106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4792_ VPWR VGND VPWR VGND uo_out[3] gpio_out_sel\[3\] net14 _1627_ _1001_ sky130_fd_sc_hd__a22o_1
XANTENNA_27 _3010_ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_38 i_tinyqv.cpu.i_core.imm_lo\[9\] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_7580_ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[23\] clknet_leaf_59_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[23\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XANTENNA_16 i_tinyqv.cpu.imm\[17\] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_6531_ VGND VPWR VPWR VGND _2943_ _2320_ _2925_ _2942_ sky130_fd_sc_hd__mux2_1
X_6462_ VPWR VGND VPWR VGND _2886_ _2885_ _2794_ _2887_ sky130_fd_sc_hd__a21o_1
X_6393_ VGND VPWR _0394_ _2831_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5413_ VPWR VGND VGND VPWR _2143_ _2128_ _1477_ sky130_fd_sc_hd__nor2_4
X_8201_ i_tinyqv.cpu.i_core.i_shift.a\[20\] clknet_leaf_40_clk _0313_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_256 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_8132_ i_tinyqv.cpu.data_addr\[7\] clknet_leaf_33_clk _0244_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_5344_ VGND VPWR _2082_ _2083_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_34_Left_115 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_8063_ i_spi.spi_dc clknet_leaf_26_clk _0198_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5275_ VGND VPWR _1313_ _2025_ _2027_ _2022_ VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4226_ VGND VPWR VPWR VGND _1073_ _1072_ i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt\[0\]
+ _1071_ sky130_fd_sc_hd__mux2_1
X_7014_ VGND VPWR VGND VPWR _3295_ _3331_ _3328_ _3304_ _3330_ _3332_ sky130_fd_sc_hd__a311o_1
XFILLER_0_49_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_4157_ VPWR VGND VGND VPWR _0985_ _1004_ _0998_ sky130_fd_sc_hd__nor2_2
Xmax_cap18 VGND VPWR _2089_ net18 VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_4088_ VPWR VGND VPWR VGND _0935_ i_tinyqv.cpu.i_core.mcause\[4\] sky130_fd_sc_hd__inv_2
X_7916_ i_tinyqv.cpu.i_core.i_registers.reg_access\[1\]\[3\] clknet_leaf_50_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[7\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7847_ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[2\] clknet_leaf_5_clk _0068_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_43_Left_124 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_65_337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_7778_ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[29\] clknet_leaf_54_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[29\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6729_ VPWR VGND VPWR VGND _3103_ _3039_ _3111_ _2995_ _1342_ _3110_ sky130_fd_sc_hd__a221o_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.i_regbuf\[23\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[23\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[27\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_191 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_52_Left_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.i_regbuf\[19\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[19\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[23\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_61_Left_142 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_70_Left_151 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.i_regbuf\[22\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[22\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[26\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_139 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_cycles.i_regbuf\[20\] i_tinyqv.cpu.i_core.i_cycles.reg_buf\[20\]
+ i_tinyqv.cpu.i_core.i_cycles.register\[24\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5060_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[5\] _1821_ _1250_ sky130_fd_sc_hd__nand2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.i_regbuf\[11\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[11\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[15\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4011_ VPWR VGND VGND VPWR _0862_ _0841_ _0861_ sky130_fd_sc_hd__or2_1
X_5962_ VGND VPWR VPWR VGND _2540_ i_tinyqv.cpu.i_core.mepc\[18\] _2504_ i_tinyqv.cpu.i_core.i_shift.a\[22\]
+ sky130_fd_sc_hd__mux2_1
X_7701_ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[16\] clknet_leaf_2_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[16\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4913_ VGND VPWR VPWR VGND _1702_ _1184_ _1701_ net198 sky130_fd_sc_hd__mux2_1
X_5893_ VGND VPWR VPWR VGND _2493_ _2492_ _2399_ i_spi.data\[4\] sky130_fd_sc_hd__mux2_1
XFILLER_0_59_186 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7632_ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[11\] clknet_leaf_44_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[11\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4844_ VGND VPWR _0036_ _1662_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_434 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7563_ i_tinyqv.cpu.i_core.i_registers.reg_access\[14\]\[2\] clknet_leaf_53_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[6\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4775_ VPWR VGND VPWR VGND _1349_ i_tinyqv.cpu.i_core.mcause\[3\] _0947_ _1610_ i_tinyqv.cpu.i_core.mstatus_mie
+ sky130_fd_sc_hd__a22o_1
X_6514_ VGND VPWR VPWR VGND _2927_ i_tinyqv.cpu.data_out\[17\] _2912_ i_tinyqv.cpu.data_out\[25\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_521 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_7494_ VPWR VGND VGND VPWR i_tinyqv.cpu.instr_data_start\[23\] _3726_ _3732_ sky130_fd_sc_hd__nor2_1
X_6445_ VGND VPWR _2825_ _2787_ _2875_ _2801_ VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_226 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_6376_ VGND VPWR VPWR VGND _2816_ i_tinyqv.mem.q_ctrl.delay_cycles_cfg\[1\] _2783_
+ _2815_ sky130_fd_sc_hd__mux2_1
X_8115_ i_tinyqv.cpu.instr_data\[0\]\[15\] clknet_leaf_12_clk _0227_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5327_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.mstatus_mte _2054_ _2070_ sky130_fd_sc_hd__nor2_1
X_8046_ i_debug_uart_tx.cycle_counter\[0\] clknet_leaf_30_clk _0181_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5258_ VPWR VGND VPWR VGND _1984_ _1981_ _2010_ _2011_ sky130_fd_sc_hd__a21o_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.i_regbuf\[8\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[8\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[12\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5189_ VPWR VGND VPWR VGND _1945_ _1944_ sky130_fd_sc_hd__inv_2
X_4209_ VGND VPWR VPWR VGND _1056_ _1055_ i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt\[1\]
+ _1053_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_0_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_5_Left_86 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_57_613 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_4_415 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4560_ VGND VPWR _1396_ _1393_ _0858_ _1395_ VPWR VGND sky130_fd_sc_hd__and3_1
X_4491_ VGND VPWR VGND VPWR _1329_ _1125_ _0846_ _1322_ _1323_ _1330_ sky130_fd_sc_hd__a311o_1
X_6230_ _2710_ _2708_ _2709_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_6161_ VGND VPWR VPWR VGND _2661_ net232 _2656_ i_tinyqv.cpu.i_core.mepc\[4\] sky130_fd_sc_hd__mux2_1
X_5112_ VPWR VGND VGND VPWR _1868_ _1871_ _1870_ sky130_fd_sc_hd__nand2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.i_regbuf\[12\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[12\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[16\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6092_ VGND VPWR VPWR VGND _2614_ i_tinyqv.cpu.i_core.i_shift.a\[18\] _2595_ i_tinyqv.cpu.i_core.i_shift.a\[22\]
+ sky130_fd_sc_hd__mux2_1
X_5043_ VPWR VGND VGND VPWR _1805_ _1803_ _1804_ sky130_fd_sc_hd__or2_1
X_6994_ VGND VPWR VGND VPWR _3314_ _3305_ _3315_ sky130_fd_sc_hd__or2_4
X_5945_ VGND VPWR VPWR VGND _2529_ _2528_ _2524_ i_tinyqv.cpu.data_addr\[12\] sky130_fd_sc_hd__mux2_1
XFILLER_0_48_613 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5876_ VGND VPWR _0226_ _2482_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4827_ VGND VPWR _0045_ _1652_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7615_ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[26\] clknet_leaf_2_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[26\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4758_ VPWR VGND VGND VPWR _1593_ _0891_ _1592_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_297 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7546_ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[21\] clknet_leaf_54_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[21\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7477_ VPWR VGND VGND VPWR i_tinyqv.cpu.data_addr\[20\] _2682_ _3005_ _3718_ sky130_fd_sc_hd__o21a_1
X_4689_ VGND VPWR VPWR VGND _1525_ _0749_ _1521_ net60 _1524_ sky130_fd_sc_hd__o2bb2a_1
X_6428_ VGND VPWR _2861_ _2860_ _2785_ _2803_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_3_481 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xi_tinyqv.cpu.i_core.i_instrret.i_regbuf\[6\] i_tinyqv.cpu.i_core.i_instrret.reg_buf\[6\]
+ i_tinyqv.cpu.i_core.i_instrret.register\[10\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6359_ VPWR VGND VGND VPWR _2800_ _1706_ _1707_ sky130_fd_sc_hd__nand2_2
XFILLER_0_11_281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_8029_ i_tinyqv.cpu.instr_data\[3\]\[7\] clknet_leaf_10_clk _0164_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_54_605 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_34_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_55_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_3991_ VPWR VGND VPWR VGND _0842_ i_tinyqv.cpu.i_core.cycle\[0\] sky130_fd_sc_hd__inv_2
X_5730_ VPWR VGND _2376_ _2333_ i_debug_uart_tx.fsm_state\[0\] i_debug_uart_tx.fsm_state\[1\]
+ i_debug_uart_tx.fsm_state\[2\] VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_29_178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_7400_ VPWR VGND VPWR VGND _3017_ _3088_ _3653_ _3650_ _3652_ _2878_ sky130_fd_sc_hd__a221o_1
X_5661_ VGND VPWR VPWR VGND _2325_ _1717_ _2308_ net272 sky130_fd_sc_hd__mux2_1
X_5592_ VGND VPWR VPWR VGND _2274_ _2275_ _2273_ _2276_ sky130_fd_sc_hd__or3_2
X_8380_ i_debug_uart_tx.uart_tx_data\[5\] clknet_leaf_19_clk _0478_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
X_4612_ VPWR VGND VPWR VGND _1447_ _1445_ _1446_ _1448_ _1408_ sky130_fd_sc_hd__a22o_1
X_4543_ VGND VPWR VPWR VGND _1381_ i_tinyqv.cpu.debug_rd\[2\] _1190_ net104 sky130_fd_sc_hd__mux2_1
X_7331_ VGND VPWR VPWR VGND _3599_ _3598_ _2147_ _3597_ sky130_fd_sc_hd__mux2_1
X_7262_ VPWR VGND VGND VPWR _2131_ _3541_ _3287_ _3535_ _3539_ _3542_ sky130_fd_sc_hd__a311o_2
X_6213_ VPWR VGND VGND VPWR _0977_ _2693_ net94 _0352_ sky130_fd_sc_hd__o21a_1
X_4474_ VPWR VGND VPWR VGND _1313_ _0842_ _1312_ sky130_fd_sc_hd__or2_2
X_7193_ VGND VPWR VGND VPWR _3490_ i_tinyqv.cpu.instr_data\[2\]\[0\] _1432_ _1418_
+ _3489_ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_473 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6144_ VGND VPWR VPWR VGND _2650_ net16 _2642_ _0814_ sky130_fd_sc_hd__mux2_1
X_6075_ VGND VPWR _0302_ _2605_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5026_ VPWR VGND VGND VPWR _1788_ _1778_ _1779_ sky130_fd_sc_hd__or2_1
X_6977_ VPWR VGND _3299_ _3298_ VPWR VGND sky130_fd_sc_hd__buf_2
X_5928_ VGND VPWR VPWR VGND _2517_ i_tinyqv.cpu.i_core.mepc\[7\] _2107_ i_tinyqv.cpu.i_core.i_shift.a\[11\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_616 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5859_ VGND VPWR VPWR VGND _2474_ i_tinyqv.cpu.instr_data\[0\]\[6\] _2469_ i_tinyqv.cpu.instr_data_in\[6\]
+ sky130_fd_sc_hd__mux2_1
X_7529_ i_tinyqv.cpu.i_core.i_registers.reg_access\[15\]\[0\] clknet_leaf_45_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[4\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.i_regbuf\[12\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[12\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[16\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_22_343 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_22_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_4190_ VGND VPWR _1036_ _1037_ _0688_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_6900_ VGND VPWR VPWR VGND _3258_ _3257_ _3254_ i_debug_uart_tx.uart_tx_data\[2\]
+ sky130_fd_sc_hd__mux2_1
X_7880_ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[3\] clknet_leaf_48_clk _0065_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_6831_ VPWR VGND VPWR VGND _3203_ _3201_ _3029_ _3204_ sky130_fd_sc_hd__a21o_1
X_6762_ VGND VPWR _3140_ _3141_ _3138_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_8501_ i_tinyqv.cpu.i_core.i_instrret.data\[3\] clknet_leaf_44_clk i_tinyqv.cpu.i_core.i_instrret.reg_buf\[7\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_3974_ VPWR VGND VPWR VGND _0821_ _0701_ _0825_ _0826_ sky130_fd_sc_hd__a21o_1
X_5713_ VPWR VGND VGND VPWR _2363_ i_debug_uart_tx.cycle_counter\[3\] _2360_ sky130_fd_sc_hd__or2_1
X_6693_ VPWR VGND VGND VPWR _3076_ _3078_ _3077_ sky130_fd_sc_hd__nand2_1
X_8432_ i_tinyqv.cpu.i_core.imm_lo\[10\] clknet_leaf_8_clk _0530_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_2
X_5644_ VGND VPWR _0163_ _2314_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8363_ i_tinyqv.cpu.instr_data_start\[21\] clknet_leaf_36_clk _0462_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_79_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5575_ VPWR VGND VGND VPWR _2266_ i_uart_rx.recieved_data\[1\] _2264_ sky130_fd_sc_hd__or2_1
Xhold211 net240 i_uart_rx.recieved_data\[6\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold200 net229 i_tinyqv.mem.qspi_data_buf\[11\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_598 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_7314_ VPWR VGND VGND VPWR net324 _3474_ _3584_ _0562_ sky130_fd_sc_hd__o21a_1
X_8294_ i_tinyqv.mem.q_ctrl.read_cycles_count\[1\] clknet_leaf_15_clk _0393_ VPWR
+ VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4526_ VPWR VGND VPWR VGND i_spi.data\[6\] _1000_ _1365_ _0997_ i_uart_rx.recieved_data\[6\]
+ _0908_ sky130_fd_sc_hd__a221o_1
Xhold244 net273 i_debug_uart_tx.uart_tx_data\[7\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold222 net251 _2085_ VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 net262 i_tinyqv.cpu.i_core.mstatus_mpie VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 net306 i_uart_rx.cycle_counter\[5\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 net295 i_tinyqv.cpu.i_core.imm_lo\[7\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4457_ VPWR VGND VGND VPWR _1030_ _1300_ _1299_ sky130_fd_sc_hd__nand2_1
Xhold255 net284 i_tinyqv.cpu.imm\[30\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7245_ VGND VPWR VPWR VGND _3528_ _3527_ _3395_ net284 sky130_fd_sc_hd__mux2_1
Xhold288 net317 i_tinyqv.mem.q_ctrl.addr\[10\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7176_ VGND VPWR VPWR VGND _3477_ _3476_ _3299_ _3328_ _3331_ _1460_ sky130_fd_sc_hd__a32o_1
X_4388_ VPWR VGND VPWR VGND _1001_ net7 _0986_ _1231_ uo_out[5] sky130_fd_sc_hd__a22o_1
X_6127_ VGND VPWR VPWR VGND _2637_ _2636_ _2468_ i_tinyqv.cpu.instr_data_in\[0\] sky130_fd_sc_hd__mux2_1
X_6058_ VGND VPWR VPWR VGND _2597_ i_tinyqv.cpu.i_core.i_shift.a\[1\] _2596_ i_tinyqv.cpu.i_core.i_shift.a\[5\]
+ sky130_fd_sc_hd__mux2_1
X_5009_ VPWR VGND VGND VPWR _1571_ _1772_ _1572_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_36_38 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_56_clk VGND VPWR clknet_3_1__leaf_clk clknet_leaf_56_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_0_42_416 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_2_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_5360_ VPWR VGND VPWR VGND _2087_ net222 _0840_ _0098_ _2095_ sky130_fd_sc_hd__a22o_1
X_5291_ VPWR VGND _2043_ _2042_ _2041_ VPWR VGND sky130_fd_sc_hd__and2_1
X_4311_ VGND VPWR VPWR VGND _1158_ _1113_ _1050_ _1111_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_368 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4242_ VGND VPWR VPWR VGND _1089_ _1087_ _1088_ _1084_ sky130_fd_sc_hd__mux2_1
X_7030_ VPWR VGND VGND VPWR _1479_ _3345_ _3282_ sky130_fd_sc_hd__nand2_1
X_4173_ VPWR VGND VGND VPWR _0957_ _1010_ _0982_ _1019_ _1020_ sky130_fd_sc_hd__o22a_1
X_7932_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[23\] clknet_leaf_36_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[23\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_47_clk VGND VPWR clknet_3_4__leaf_clk clknet_leaf_47_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_7863_ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[18\] clknet_leaf_3_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[18\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6814_ VPWR VGND VGND VPWR _0784_ _3188_ i_tinyqv.cpu.imm\[18\] sky130_fd_sc_hd__nand2_1
X_7794_ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[13\] clknet_leaf_57_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[13\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6745_ _3125_ _3116_ _3105_ _3117_ _3114_ VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_0_45_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_3957_ VPWR VGND VPWR VGND _0690_ i_tinyqv.cpu.imm\[22\] _0619_ _0809_ i_tinyqv.cpu.imm\[26\]
+ sky130_fd_sc_hd__a22o_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.i_regbuf\[26\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[26\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[30\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6676_ VPWR VGND VPWR VGND _3062_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[14\]
+ sky130_fd_sc_hd__inv_2
X_3888_ VGND VPWR VGND VPWR i_tinyqv.cpu.i_core.i_registers.reg_access\[1\]\[0\] _0740_
+ _0739_ _0738_ _0648_ _0737_ sky130_fd_sc_hd__a2111oi_4
X_8415_ i_tinyqv.cpu.is_store clknet_leaf_7_clk _0513_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_5627_ VPWR VGND VPWR VGND i_tinyqv.mem.q_ctrl.is_writing _2302_ _1543_ _2303_ sky130_fd_sc_hd__a21o_1
X_5558_ VPWR VGND VGND VPWR _2253_ _2254_ _0137_ sky130_fd_sc_hd__nor2_1
X_8346_ i_tinyqv.cpu.instr_data_start\[4\] clknet_leaf_24_clk _0445_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
X_8277_ i_tinyqv.mem.data_from_read\[17\] clknet_leaf_13_clk _0376_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_4509_ VPWR VGND VPWR VGND _1348_ _0933_ _0930_ sky130_fd_sc_hd__or2_2
X_5489_ _2203_ _2200_ _2205_ _2204_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.i_regbuf\[15\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[15\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[19\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7228_ VPWR VGND _3517_ _3408_ _3330_ _3328_ _3510_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_7159_ VGND VPWR VPWR VGND _3462_ _3461_ _3396_ i_tinyqv.cpu.i_core.imm_lo\[10\]
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_38_clk VGND VPWR clknet_3_4__leaf_clk clknet_leaf_38_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_64_541 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_32_460 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_29_clk VGND VPWR clknet_3_7__leaf_clk clknet_leaf_29_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_4860_ VGND VPWR _0079_ _1671_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_3811_ VPWR VGND _0663_ i_tinyqv.cpu.i_core.i_registers.rs2\[1\] VPWR VGND sky130_fd_sc_hd__buf_6
XANTENNA_28 i_debug_uart_tx.uart_tx_data\[2\] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_6530_ VGND VPWR VPWR VGND _2942_ _2941_ _2792_ _2939_ sky130_fd_sc_hd__mux2_1
X_4791_ VPWR VGND VPWR VGND _1012_ i_tinyqv.cpu.instr_data_in\[3\] _1625_ _1626_ sky130_fd_sc_hd__a21o_1
XANTENNA_39 i_tinyqv.cpu.i_core.imm_lo\[9\] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_17 i_tinyqv.cpu.imm\[20\] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_6461_ VGND VPWR VPWR VGND _2886_ _2836_ _2803_ _1715_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_544 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_70_533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_15_449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_6392_ VGND VPWR VPWR VGND _2831_ _2830_ _2811_ i_tinyqv.mem.q_ctrl.read_cycles_count\[2\]
+ sky130_fd_sc_hd__mux2_1
X_8200_ i_tinyqv.cpu.i_core.i_shift.a\[19\] clknet_leaf_40_clk _0312_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5412_ VPWR VGND VGND VPWR _1490_ _1507_ _2142_ sky130_fd_sc_hd__nor2_1
X_8131_ i_tinyqv.cpu.data_addr\[6\] clknet_leaf_32_clk _0243_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_5343_ VPWR VGND VPWR VGND i_tinyqv.cpu.i_core.is_double_fault_r _2070_ _1400_ _2082_
+ sky130_fd_sc_hd__or3_1
X_8062_ i_spi.busy clknet_leaf_27_clk _0197_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5274_ VPWR VGND VPWR VGND _1313_ _2025_ _2022_ _2026_ sky130_fd_sc_hd__or3_1
X_4225_ VGND VPWR VPWR VGND _1072_ i_tinyqv.cpu.i_core.i_shift.a\[23\] _1027_ i_tinyqv.cpu.i_core.i_shift.a\[8\]
+ sky130_fd_sc_hd__mux2_1
X_7013_ VGND VPWR VPWR VGND _3308_ _3331_ _2126_ sky130_fd_sc_hd__and2b_2
X_4156_ VPWR VGND VGND VPWR _0983_ _0995_ _0984_ _1003_ sky130_fd_sc_hd__nor3_1
Xmax_cap19 VGND VPWR net19 _0948_ VPWR VGND sky130_fd_sc_hd__buf_1
X_4087_ VPWR VGND VGND VPWR _0934_ _0933_ _0922_ sky130_fd_sc_hd__or2_1
X_7915_ i_tinyqv.cpu.i_core.i_registers.reg_access\[1\]\[2\] clknet_leaf_50_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[6\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7846_ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[1\] clknet_leaf_5_clk _0067_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.i_regbuf\[27\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[27\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[31\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7777_ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[28\] clknet_leaf_0_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[28\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4989_ VPWR VGND _1753_ _1752_ VPWR VGND sky130_fd_sc_hd__buf_4
XFILLER_0_46_552 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_6728_ VGND VPWR VGND VPWR _3110_ _3040_ _3108_ _3109_ _3047_ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_298 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_6659_ VGND VPWR net40 _3047_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_8329_ i_tinyqv.mem.q_ctrl.last_ram_a_sel clknet_leaf_17_clk _0428_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.i_regbuf\[16\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[16\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[20\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.i_regbuf\[30\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[30\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[2\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_107 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_24_246 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.i_regbuf\[15\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[15\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[19\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_485 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xi_tinyqv.cpu.i_core.i_cycles.i_regbuf\[13\] i_tinyqv.cpu.i_core.i_cycles.reg_buf\[13\]
+ i_tinyqv.cpu.i_core.i_cycles.register\[17\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4010_ VGND VPWR VGND VPWR _0860_ _0848_ _0850_ _0861_ sky130_fd_sc_hd__o21ba_1
X_5961_ VGND VPWR _0254_ _2539_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7700_ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[15\] clknet_leaf_58_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[15\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4912_ _1647_ _1701_ _1188_ _1695_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_47_305 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5892_ VGND VPWR VPWR VGND _2492_ i_spi.data\[3\] _2386_ i_debug_uart_tx.uart_tx_data\[4\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7631_ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[10\] clknet_leaf_45_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[10\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4843_ VGND VPWR VPWR VGND _1662_ i_tinyqv.cpu.debug_rd\[2\] _1659_ i_tinyqv.cpu.i_core.i_registers.reg_access\[11\]\[2\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_179 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7562_ i_tinyqv.cpu.i_core.i_registers.reg_access\[14\]\[1\] clknet_leaf_57_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[5\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_202 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4774_ VPWR VGND VGND VPWR _0939_ _1348_ _1609_ sky130_fd_sc_hd__nor2_1
X_6513_ VGND VPWR _0419_ _2926_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7493_ VPWR VGND VPWR VGND _3730_ i_tinyqv.mem.q_ctrl.addr\[22\] _3009_ _0594_ _3731_
+ sky130_fd_sc_hd__a22o_1
X_6444_ VGND VPWR _0402_ _2874_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_9_clk VGND VPWR clknet_3_2__leaf_clk clknet_leaf_9_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_6375_ VGND VPWR VGND VPWR i_tinyqv.mem.q_ctrl.read_cycles_count\[1\] _2796_ _2815_
+ _2814_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_11_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_3_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_8114_ i_tinyqv.cpu.instr_data\[0\]\[14\] clknet_leaf_12_clk _0226_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5326_ VPWR VGND VPWR VGND _2069_ _2064_ _2067_ _0090_ sky130_fd_sc_hd__a21oi_1
X_8045_ i_debug_uart_tx.data_to_send\[7\] clknet_leaf_28_clk _0180_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5257_ VPWR VGND VGND VPWR _2008_ _2010_ _2009_ sky130_fd_sc_hd__nand2_1
X_4208_ VGND VPWR VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[24\] i_tinyqv.cpu.i_core.i_shift.a\[25\]
+ i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt\[0\] _1054_ i_tinyqv.cpu.i_core.i_shift.a\[6\]
+ _1029_ _1055_ sky130_fd_sc_hd__mux4_1
X_5188_ VPWR VGND _1944_ _1943_ _1942_ VPWR VGND sky130_fd_sc_hd__and2_1
X_4139_ VPWR VGND VGND VPWR _0985_ _0986_ _0983_ sky130_fd_sc_hd__nor2_2
X_7829_ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[16\] clknet_leaf_49_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[16\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.i_regbuf\[31\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[31\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[3\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.i_regbuf\[20\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[20\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[24\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.i_regbuf\[27\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[27\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[31\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_647 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xclkbuf_3_4__f_clk VGND VPWR VGND VPWR clknet_0_clk clknet_3_4__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_72_628 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_56_157 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_37_393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_4490_ VPWR VGND VPWR VGND _1328_ _1326_ _0847_ _1329_ sky130_fd_sc_hd__a21oi_1
X_6160_ VGND VPWR _0332_ _2660_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5111_ VGND VPWR _1846_ _1869_ _1870_ _1844_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_6091_ VGND VPWR _0310_ _2613_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5042_ VPWR VGND VPWR VGND _1788_ _1776_ _1802_ _1804_ sky130_fd_sc_hd__a21oi_1
X_6993_ VGND VPWR VPWR VGND _3313_ _1465_ _2155_ _3314_ sky130_fd_sc_hd__or3_2
X_5944_ VGND VPWR VPWR VGND _2528_ i_tinyqv.cpu.i_core.mepc\[12\] _2504_ i_tinyqv.cpu.i_core.i_shift.a\[16\]
+ sky130_fd_sc_hd__mux2_1
X_5875_ VGND VPWR VPWR VGND _2482_ net266 _2468_ _1720_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_146 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7614_ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[25\] clknet_leaf_52_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[25\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4826_ VGND VPWR VPWR VGND _1652_ i_tinyqv.cpu.debug_rd\[3\] _1648_ i_tinyqv.cpu.i_core.i_registers.reg_access\[13\]\[3\]
+ sky130_fd_sc_hd__mux2_1
X_7545_ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[20\] clknet_leaf_47_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[20\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4757_ VPWR VGND VPWR VGND _0890_ _0883_ i_tinyqv.cpu.instr_data_start\[7\] _1592_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_276 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4688_ VPWR VGND VGND VPWR _1522_ _1524_ _1523_ sky130_fd_sc_hd__nand2_1
X_7476_ VPWR VGND VPWR VGND _3017_ _3211_ _3717_ _3714_ _3716_ _2878_ sky130_fd_sc_hd__a221o_1
X_6427_ VPWR VGND VPWR VGND _2860_ _2794_ sky130_fd_sc_hd__inv_2
X_6358_ VPWR VGND VPWR VGND _2794_ _2798_ _2795_ _2790_ _2799_ sky130_fd_sc_hd__or4_1
X_5309_ VGND VPWR VGND VPWR _1392_ _1394_ i_tinyqv.cpu.i_core.is_interrupt _2056_
+ sky130_fd_sc_hd__a21o_2
X_6289_ VGND VPWR VPWR VGND _2754_ _2318_ _1552_ i_tinyqv.mem.qspi_data_buf\[9\] sky130_fd_sc_hd__mux2_1
X_8028_ i_tinyqv.cpu.instr_data\[3\]\[6\] clknet_leaf_4_clk _0163_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_625 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_38_135 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_30_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.i_regbuf\[5\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[5\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[9\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3990_ VPWR VGND VGND VPWR _0841_ _0838_ _0840_ sky130_fd_sc_hd__nand2_2
X_5660_ VGND VPWR _0169_ _2324_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_4611_ VGND VPWR VPWR VGND _1447_ i_tinyqv.cpu.instr_data\[2\]\[3\] _1412_ i_tinyqv.cpu.instr_data\[0\]\[3\]
+ sky130_fd_sc_hd__mux2_1
X_5591_ VPWR VGND VPWR VGND i_uart_rx.cycle_counter\[5\] i_uart_rx.cycle_counter\[3\]
+ _2275_ i_uart_rx.cycle_counter\[2\] i_uart_rx.cycle_counter\[4\] sky130_fd_sc_hd__or4bb_1
X_4542_ VPWR VGND i_tinyqv.cpu.debug_rd\[2\] _1380_ VPWR VGND sky130_fd_sc_hd__buf_4
X_7330_ VGND VPWR VPWR VGND _3598_ _3556_ _3454_ _1491_ _3390_ _3290_ sky130_fd_sc_hd__a32o_1
X_4473_ VPWR VGND net44 _1312_ net65 VPWR VGND sky130_fd_sc_hd__and2_2
X_7261_ _3541_ _2123_ _3335_ _3532_ _3540_ _3531_ VPWR VGND VGND VPWR sky130_fd_sc_hd__o311a_1
X_6212_ VPWR VGND VPWR VGND _2692_ i_tinyqv.mem.data_stall _2691_ _2693_ i_tinyqv.mem.q_ctrl.data_req
+ sky130_fd_sc_hd__a22o_1
X_7192_ VPWR VGND VGND VPWR _3487_ _3488_ _3489_ sky130_fd_sc_hd__nor2_1
X_6143_ VGND VPWR _0326_ _2649_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6074_ VGND VPWR VPWR VGND _2605_ i_tinyqv.cpu.i_core.i_shift.a\[13\] _2593_ i_tinyqv.cpu.i_core.i_shift.a\[9\]
+ sky130_fd_sc_hd__mux2_1
X_5025_ VPWR VGND VPWR VGND _1785_ _1783_ _1786_ _1787_ sky130_fd_sc_hd__a21o_1
X_6976_ VPWR VGND VPWR VGND _1503_ _1461_ _1506_ _3298_ sky130_fd_sc_hd__a21o_1
X_5927_ VGND VPWR _0243_ _2516_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_433 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_8_541 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5858_ VGND VPWR _0217_ _2473_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5789_ VPWR VGND VPWR VGND _2398_ i_spi.spi_clk_out _2395_ _2423_ _2403_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_585 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Right_17 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4809_ VPWR VGND _1189_ _1642_ _1641_ VPWR VGND sky130_fd_sc_hd__and2_2
X_7528_ VPWR VGND VPWR VGND _3746_ net90 _3754_ _0606_ sky130_fd_sc_hd__a21oi_1
X_7459_ VGND VPWR _3697_ _3702_ _0784_ VPWR VGND sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_26_Right_26 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xsplit31 VGND VPWR net60 i_tinyqv.cpu.pc\[2\] VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_35_Right_35 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_54_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_44_Right_44 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6830_ VGND VPWR VGND VPWR _3203_ _2987_ _3202_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[27\]
+ _2993_ sky130_fd_sc_hd__a211o_1
X_6761_ VPWR VGND VGND VPWR _3126_ _3139_ _3140_ sky130_fd_sc_hd__nor2_1
X_5712_ VGND VPWR _0183_ _2362_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_53_Right_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_8500_ i_tinyqv.cpu.i_core.i_instrret.data\[2\] clknet_leaf_49_clk i_tinyqv.cpu.i_core.i_instrret.reg_buf\[6\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_3973_ VPWR VGND VPWR VGND _0824_ _0656_ net141 _0825_ sky130_fd_sc_hd__a21oi_1
X_6692_ VPWR VGND VGND VPWR _3077_ i_tinyqv.cpu.instr_data_start\[7\] i_tinyqv.cpu.i_core.imm_lo\[7\]
+ sky130_fd_sc_hd__or2_1
X_8431_ VGND VPWR VGND VPWR i_tinyqv.cpu.i_core.imm_lo\[9\] _0529_ clknet_leaf_8_clk
+ sky130_fd_sc_hd__dfxtp_4
X_5643_ VGND VPWR VPWR VGND _2314_ i_tinyqv.cpu.instr_data_in\[6\] _2309_ i_tinyqv.cpu.instr_data\[3\]\[6\]
+ sky130_fd_sc_hd__mux2_1
X_5574_ VGND VPWR VGND VPWR _0142_ net201 _2263_ _2265_ _2240_ sky130_fd_sc_hd__o211a_1
X_8362_ i_tinyqv.cpu.instr_data_start\[20\] clknet_leaf_36_clk _0461_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
X_4525_ VPWR VGND VPWR VGND net8 _0986_ _1364_ net14 gpio_out_sel\[6\] _1363_ sky130_fd_sc_hd__a221o_1
X_7313_ VPWR VGND VPWR VGND _3504_ _3583_ _3362_ _3584_ sky130_fd_sc_hd__or3_1
Xhold201 net230 i_tinyqv.cpu.i_core.mie\[16\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_8293_ i_tinyqv.mem.q_ctrl.read_cycles_count\[0\] clknet_leaf_15_clk _0392_ VPWR
+ VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
Xhold212 net241 i_uart_rx.recieved_data\[3\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 net263 i_tinyqv.cpu.instr_data\[3\]\[2\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 net252 i_tinyqv.cpu.i_core.i_registers.rd\[3\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 net274 i_tinyqv.mem.q_ctrl.spi_in_buffer\[7\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 net307 i_uart_rx.cycle_counter\[1\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold256 net285 i_tinyqv.mem.data_from_read\[23\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4456_ VPWR VGND _1299_ _1298_ _1289_ _1046_ _1121_ VGND VPWR sky130_fd_sc_hd__a31o_1
Xhold267 net296 i_tinyqv.cpu.i_core.imm_lo\[11\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7244_ VPWR VGND _3527_ _3460_ _3330_ _3291_ _3509_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_4387_ VPWR VGND VPWR VGND i_spi.data\[1\] _1000_ _1230_ _0986_ net3 _1229_ sky130_fd_sc_hd__a221o_1
Xhold289 net318 i_tinyqv.mem.q_ctrl.addr\[15\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7175_ VPWR VGND VGND VPWR _3476_ _1467_ _3315_ sky130_fd_sc_hd__nand2_2
X_6126_ VPWR VGND VGND VPWR _2636_ _1400_ i_tinyqv.cpu.instr_data\[0\]\[0\] sky130_fd_sc_hd__or2_1
X_6057_ VGND VPWR _2595_ _2596_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_5008_ VGND VPWR _1770_ _1771_ _1769_ VPWR VGND sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_71_Right_71 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6959_ VGND VPWR _3281_ _3282_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_23_108 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_80_Right_80 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_35_491 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_2_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_22_152 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_77_24 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_50_472 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5290_ VPWR VGND VGND VPWR _2042_ _2039_ _2040_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_4310_ VGND VPWR VPWR VGND _1157_ _1110_ _1050_ _1106_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4241_ VGND VPWR i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt\[1\] _1088_ VPWR
+ VGND sky130_fd_sc_hd__clkbuf_4
X_4172_ VGND VPWR VPWR VGND _1019_ _1018_ _0907_ _1013_ sky130_fd_sc_hd__mux2_1
X_7931_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[22\] clknet_leaf_36_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[22\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_50 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7862_ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[17\] clknet_leaf_47_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[17\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6813_ VPWR VGND VGND VPWR _0784_ i_tinyqv.cpu.imm\[18\] _3187_ sky130_fd_sc_hd__nor2_1
X_7793_ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[12\] clknet_leaf_2_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[12\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_583 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_58_572 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_18_414 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_3956_ VPWR VGND VGND VPWR _0807_ _0803_ _0801_ _0808_ sky130_fd_sc_hd__nor3_1
X_6744_ VPWR VGND VPWR VGND _3124_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[20\]
+ sky130_fd_sc_hd__inv_2
X_6675_ VGND VPWR VGND VPWR _0446_ i_tinyqv.cpu.instr_data_start\[5\] _3027_ _3061_
+ _2061_ sky130_fd_sc_hd__o211a_1
X_5626_ VPWR VGND VPWR VGND _2302_ i_tinyqv.mem.q_ctrl.spi_clk_out sky130_fd_sc_hd__inv_2
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.i_regbuf\[19\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[19\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[23\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_330 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_3887_ VPWR VGND VPWR VGND _0638_ i_tinyqv.cpu.i_core.i_registers.reg_access\[8\]\[0\]
+ net321 _0739_ i_tinyqv.cpu.i_core.i_registers.reg_access\[2\]\[0\] sky130_fd_sc_hd__a22o_1
X_8414_ i_tinyqv.cpu.is_auipc clknet_leaf_6_clk _0512_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5557_ VGND VPWR _2251_ _2242_ _2254_ i_uart_rx.cycle_counter\[6\] VPWR VGND sky130_fd_sc_hd__o21ai_1
X_8345_ i_tinyqv.cpu.instr_data_start\[3\] clknet_leaf_24_clk _0444_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5488_ VPWR VGND _2204_ _2197_ i_uart_tx.cycle_counter\[0\] net206 i_uart_tx.cycle_counter\[2\]
+ VGND VPWR sky130_fd_sc_hd__a31o_1
X_8276_ i_tinyqv.mem.data_from_read\[16\] clknet_leaf_13_clk _0375_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_697 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4508_ VPWR VGND VPWR VGND _1346_ _1336_ _0858_ _1347_ sky130_fd_sc_hd__a21o_1
X_4439_ VGND VPWR VPWR VGND _1282_ _1134_ _1108_ _1281_ sky130_fd_sc_hd__mux2_1
X_7227_ VPWR VGND VPWR VGND _3515_ _3474_ _3516_ _0543_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_71 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7158_ VPWR VGND VPWR VGND _1478_ _1514_ _3461_ _3364_ _3460_ _3456_ sky130_fd_sc_hd__a221o_1
X_6109_ VGND VPWR _0319_ _2622_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7089_ VPWR VGND VPWR VGND _2130_ _2133_ _2121_ _3399_ sky130_fd_sc_hd__or3_1
XFILLER_0_49_583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_2_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_4790_ VPWR VGND _1625_ _0979_ _0869_ i_tinyqv.cpu.instr_data_in\[11\] _0865_ VGND
+ VPWR sky130_fd_sc_hd__a31o_1
X_3810_ VPWR VGND _0662_ i_tinyqv.cpu.i_core.i_registers.rs2\[0\] VPWR VGND sky130_fd_sc_hd__buf_2
XANTENNA_18 i_tinyqv.mem.q_ctrl.addr\[21\] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_29 i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[3\] VGND VPWR VPWR VGND
+ sky130_fd_sc_hd__diode_2
X_6460_ VGND VPWR VGND VPWR _2885_ _2884_ _2803_ _2800_ _2813_ sky130_fd_sc_hd__a211o_1
XFILLER_0_12_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6391_ VGND VPWR VGND VPWR _2823_ _2827_ _2828_ _2830_ _2829_ sky130_fd_sc_hd__a2bb2o_1
X_5411_ VGND VPWR VGND VPWR _2141_ _1469_ _2124_ _2139_ _2140_ sky130_fd_sc_hd__o211a_1
X_5342_ VPWR VGND VGND VPWR _0956_ _2081_ _1619_ sky130_fd_sc_hd__nand2_1
X_8130_ i_tinyqv.cpu.data_addr\[5\] clknet_leaf_25_clk _0242_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_344 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_8061_ i_spi.bits_remaining\[3\] clknet_leaf_26_clk net195 VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5273_ VGND VPWR _2024_ _2025_ _2023_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_7012_ VPWR VGND _3330_ _3329_ VPWR VGND sky130_fd_sc_hd__buf_2
X_4224_ VGND VPWR VPWR VGND _1071_ i_tinyqv.cpu.i_core.i_shift.a\[22\] _1027_ i_tinyqv.cpu.i_core.i_shift.a\[9\]
+ sky130_fd_sc_hd__mux2_1
X_4155_ VPWR VGND VPWR VGND _1001_ i_spi.data\[0\] _1000_ _1002_ uo_out[0] sky130_fd_sc_hd__a22o_1
X_4086_ VPWR VGND VPWR VGND _0932_ _0933_ i_tinyqv.cpu.i_core.imm_lo\[6\] _0923_ sky130_fd_sc_hd__or3b_2
X_7914_ i_tinyqv.cpu.i_core.i_registers.reg_access\[1\]\[1\] clknet_leaf_51_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[5\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7845_ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[0\] clknet_leaf_48_clk _0066_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7776_ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[27\] clknet_leaf_58_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[27\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4988_ VPWR VGND _1752_ i_tinyqv.cpu.i_core.i_cycles.rstn VPWR VGND sky130_fd_sc_hd__buf_4
X_6727_ VPWR VGND VGND VPWR _1390_ _3109_ _2523_ sky130_fd_sc_hd__nand2_1
X_3939_ _0791_ _0732_ _0611_ _0690_ _0733_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
XFILLER_0_46_564 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_6658_ VPWR VGND VGND VPWR _1390_ _3046_ _2511_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_288 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5609_ VPWR VGND VGND VPWR _2290_ i_uart_rx.fsm_state\[1\] i_uart_rx.fsm_state\[0\]
+ sky130_fd_sc_hd__or2_1
X_8328_ i_tinyqv.mem.q_ctrl.last_ram_b_sel clknet_leaf_17_clk _0427_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_6589_ VGND VPWR net31 _2987_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_8259_ VGND VPWR VGND VPWR i_tinyqv.mem.qspi_data_byte_idx\[1\] _0358_ clknet_leaf_17_clk
+ sky130_fd_sc_hd__dfxtp_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.i_regbuf\[23\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[23\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[27\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_634 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_68_122 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.i_regbuf\[12\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[12\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[16\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_37_586 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_74_25 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_instrret.i_regbuf\[22\] i_tinyqv.cpu.i_core.i_instrret.reg_buf\[22\]
+ i_tinyqv.cpu.i_core.i_instrret.register\[26\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5960_ VGND VPWR VPWR VGND _2539_ _2538_ _2524_ i_tinyqv.cpu.data_addr\[17\] sky130_fd_sc_hd__mux2_1
X_5891_ VGND VPWR _0232_ _2491_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4911_ VGND VPWR _0061_ _1700_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7630_ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[9\] clknet_leaf_55_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[9\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4842_ VGND VPWR _0035_ _1661_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7561_ i_tinyqv.cpu.i_core.i_registers.reg_access\[14\]\[0\] clknet_leaf_57_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[4\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_458 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4773_ VPWR VGND VPWR VGND _1607_ i_tinyqv.cpu.i_core.cycle_count\[3\] _0931_ _1608_
+ _0927_ sky130_fd_sc_hd__a22o_1
X_7492_ VPWR VGND VPWR VGND _3007_ i_tinyqv.mem.q_ctrl.addr\[18\] _3005_ _3731_ sky130_fd_sc_hd__a21o_1
X_6512_ VGND VPWR VPWR VGND _2926_ _2316_ _2925_ _2922_ sky130_fd_sc_hd__mux2_1
X_6443_ VPWR VGND _2874_ _2873_ _2832_ VPWR VGND sky130_fd_sc_hd__and2_1
X_6374_ VPWR VGND VPWR VGND i_tinyqv.mem.q_ctrl.read_cycles_count\[2\] _2796_ i_tinyqv.mem.q_ctrl.read_cycles_count\[1\]
+ _2814_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_8113_ i_tinyqv.cpu.instr_data\[0\]\[13\] clknet_leaf_13_clk _0225_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5325_ VPWR VGND VGND VPWR net158 _2069_ _2054_ sky130_fd_sc_hd__nand2_1
X_8044_ i_debug_uart_tx.data_to_send\[6\] clknet_leaf_28_clk _0179_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5256_ VPWR VGND VGND VPWR _2009_ i_tinyqv.cpu.i_core.multiplier.accum\[14\] _2007_
+ sky130_fd_sc_hd__or2_1
X_4207_ VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[7\] _1054_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_5187_ VGND VPWR _1916_ _1913_ _1943_ _1915_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_4138_ VPWR VGND VPWR VGND _0985_ _0984_ _0969_ sky130_fd_sc_hd__or2_2
X_4069_ VPWR VGND VGND VPWR _0689_ _0916_ _0688_ sky130_fd_sc_hd__nand2_4
X_7828_ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[15\] clknet_leaf_52_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[15\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7759_ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[10\] clknet_leaf_53_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[10\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.i_regbuf\[24\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[24\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[28\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.i_regbuf\[13\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[13\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[17\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_65_681 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_25_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_5110_ VGND VPWR VGND VPWR _1841_ _1869_ _1843_ sky130_fd_sc_hd__or2b_1
X_6090_ VGND VPWR VPWR VGND _2613_ i_tinyqv.cpu.i_core.i_shift.a\[17\] _2596_ i_tinyqv.cpu.i_core.i_shift.a\[21\]
+ sky130_fd_sc_hd__mux2_1
X_5041_ VGND VPWR _1803_ _1788_ _1776_ _1802_ VPWR VGND sky130_fd_sc_hd__and3_1
X_6992_ VPWR VGND VPWR VGND _3313_ _1460_ sky130_fd_sc_hd__inv_2
X_5943_ VGND VPWR _0248_ _2527_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_103 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5874_ VGND VPWR _0225_ _2481_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_501 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7613_ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[24\] clknet_leaf_0_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[24\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4825_ VGND VPWR _0044_ _1651_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7544_ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[19\] clknet_leaf_46_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[19\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4756_ VGND VPWR VPWR VGND _0884_ _1591_ _0888_ sky130_fd_sc_hd__xor2_1
X_4687_ VPWR VGND VGND VPWR _1523_ i_tinyqv.cpu.instr_write_offset\[2\] _1519_ sky130_fd_sc_hd__or2_1
X_7475_ VPWR VGND VGND VPWR _3017_ _3715_ _3716_ sky130_fd_sc_hd__nor2_1
X_6426_ VGND VPWR _0399_ _2859_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.i_regbuf\[6\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[6\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[10\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6357_ VGND VPWR VPWR VGND _2798_ _2796_ _2797_ i_tinyqv.mem.q_ctrl.delay_cycles_cfg\[0\]
+ sky130_fd_sc_hd__mux2_1
X_5308_ VPWR VGND VGND VPWR _2055_ i_tinyqv.cpu.i_core.is_interrupt _2054_ sky130_fd_sc_hd__or2_1
X_6288_ VGND VPWR _0367_ _2753_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5239_ VPWR VGND VGND VPWR _1991_ _1993_ _1992_ sky130_fd_sc_hd__nand2_1
X_8027_ i_tinyqv.cpu.instr_data\[3\]\[5\] clknet_leaf_3_clk _0162_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_629 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_49_Left_130 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_39_28 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.i_regbuf\[5\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[5\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[9\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4610_ VPWR VGND VGND VPWR i_tinyqv.cpu.instr_data\[1\]\[3\] _1414_ _1416_ _1446_
+ sky130_fd_sc_hd__o21a_1
X_5590_ VPWR VGND VPWR VGND i_uart_rx.cycle_counter\[7\] i_uart_rx.cycle_counter\[6\]
+ i_uart_rx.cycle_counter\[1\] _2274_ i_uart_rx.cycle_counter\[0\] sky130_fd_sc_hd__or4b_1
XFILLER_0_25_353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_4541_ VGND VPWR VGND VPWR _1380_ _1332_ _1330_ _0877_ _1379_ _1034_ sky130_fd_sc_hd__a32o_2
XFILLER_0_20_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4472_ VPWR VGND VPWR VGND _1311_ i_tinyqv.cpu.i_core.i_shift.a\[2\] sky130_fd_sc_hd__inv_2
X_7260_ VPWR VGND VGND VPWR _3540_ _2124_ _3467_ sky130_fd_sc_hd__or2_1
X_6211_ VGND VPWR VPWR VGND _2692_ _0870_ _0867_ _0871_ sky130_fd_sc_hd__mux2_1
X_7191_ VPWR VGND VGND VPWR _1461_ _3488_ _1504_ sky130_fd_sc_hd__nor2_2
X_6142_ VGND VPWR VPWR VGND _2649_ _2648_ _2645_ _1149_ sky130_fd_sc_hd__mux2_1
X_6073_ VGND VPWR _0301_ _2604_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5024_ VPWR VGND _1786_ _1782_ _1780_ VPWR VGND sky130_fd_sc_hd__and2_1
X_6975_ VPWR VGND VGND VPWR _3297_ _1483_ _2127_ sky130_fd_sc_hd__or2_1
X_5926_ VGND VPWR VPWR VGND _2516_ _2515_ _2502_ i_tinyqv.cpu.data_addr\[6\] sky130_fd_sc_hd__mux2_1
X_5857_ VGND VPWR VPWR VGND _2473_ i_tinyqv.cpu.instr_data\[0\]\[5\] _2469_ i_tinyqv.cpu.instr_data_in\[5\]
+ sky130_fd_sc_hd__mux2_1
X_5788_ VPWR VGND VGND VPWR _2421_ _2418_ _0199_ _2394_ _2221_ _2422_ sky130_fd_sc_hd__o221ai_1
X_4808_ VPWR VGND _1641_ _1640_ i_tinyqv.cpu.i_core.i_registers.rd\[1\] VPWR VGND
+ sky130_fd_sc_hd__and2_1
X_4739_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[3\] _1574_ _1166_ sky130_fd_sc_hd__nand2_1
X_7527_ VGND VPWR _3746_ _2079_ _3754_ net90 VPWR VGND sky130_fd_sc_hd__o21ai_1
X_7458_ VPWR VGND VGND VPWR _3625_ net301 _3624_ net304 _0589_ _3701_ sky130_fd_sc_hd__o221a_1
XFILLER_0_16_386 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_6409_ VGND VPWR _2845_ _2792_ i_tinyqv.mem.q_ctrl.spi_flash_select _1709_ VPWR VGND
+ sky130_fd_sc_hd__and3_1
X_7389_ VPWR VGND VGND VPWR net126 _3624_ _2733_ _3644_ sky130_fd_sc_hd__o21a_1
XFILLER_0_12_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_31_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_39_401 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_35_640 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_58_710 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6760_ _3139_ _3116_ _3105_ _3117_ _3114_ _3127_ VPWR VGND VGND VPWR sky130_fd_sc_hd__o311a_1
X_5711_ _2360_ _2357_ _2362_ _2361_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_3972_ VPWR VGND VGND VPWR _0824_ _0822_ _0823_ sky130_fd_sc_hd__nand2_2
X_6691_ VPWR VGND VGND VPWR i_tinyqv.cpu.instr_data_start\[7\] _3076_ i_tinyqv.cpu.i_core.imm_lo\[7\]
+ sky130_fd_sc_hd__nand2_1
X_5642_ VGND VPWR _0162_ _2313_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8430_ i_tinyqv.cpu.i_core.imm_lo\[8\] clknet_leaf_23_clk _0528_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_2
X_5573_ VPWR VGND VGND VPWR _2265_ i_uart_rx.recieved_data\[0\] _2264_ sky130_fd_sc_hd__or2_1
X_8361_ i_tinyqv.cpu.instr_data_start\[19\] clknet_leaf_36_clk _0460_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
X_4524_ VPWR VGND _1363_ uo_out[6] _1001_ VPWR VGND sky130_fd_sc_hd__and2_1
Xhold202 net231 i_tinyqv.cpu.imm\[14\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_695 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7312_ VPWR VGND VGND VPWR _2165_ _3571_ _3572_ _3583_ sky130_fd_sc_hd__o21a_1
Xhold224 net253 i_tinyqv.mem.qspi_data_buf\[27\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_8292_ i_tinyqv.cpu.instr_fetch_started clknet_leaf_20_clk _0391_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_367 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold213 net242 i_tinyqv.cpu.additional_mem_ops\[1\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 net264 i_tinyqv.cpu.i_core.mepc\[5\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 net286 i_tinyqv.mem.qspi_data_buf\[25\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 net275 i_tinyqv.mem.qspi_data_buf\[8\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 net297 i_tinyqv.cpu.data_addr\[7\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4455_ VGND VPWR VGND VPWR _1048_ _1297_ _1077_ _1291_ _1293_ _1298_ sky130_fd_sc_hd__a311o_1
X_7243_ VPWR VGND VGND VPWR net146 _3360_ _3526_ _0549_ sky130_fd_sc_hd__o21a_1
X_4386_ VGND VPWR VPWR VGND _1229_ _1228_ _0987_ _1225_ _1003_ gpio_out_sel\[1\] sky130_fd_sc_hd__a32o_1
Xhold279 net308 i_spi.end_txn_reg VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7174_ VGND VPWR VGND VPWR _3475_ _3465_ _3472_ _3364_ _3362_ sky130_fd_sc_hd__a211o_1
X_6125_ VGND VPWR _0322_ _2635_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6056_ VGND VPWR VGND VPWR _1563_ _1031_ _2595_ _1124_ sky130_fd_sc_hd__a21oi_4
X_5007_ VPWR VGND _1770_ _1166_ i_tinyqv.cpu.i_core.i_shift.a\[4\] VPWR VGND sky130_fd_sc_hd__and2_1
X_6958_ VPWR VGND _3281_ _3280_ VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_0_48_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6889_ VGND VPWR VGND VPWR _3251_ net294 _0957_ i_tinyqv.cpu.data_write_n\[1\] _0979_
+ sky130_fd_sc_hd__a211o_1
X_5909_ VGND VPWR _2106_ _2504_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_8559_ i_tinyqv.cpu.i_core.i_shift.b\[4\] clknet_leaf_40_clk _0601_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_6_309 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4240_ VGND VPWR VPWR VGND _1087_ _1086_ _1083_ _1085_ sky130_fd_sc_hd__mux2_1
X_4171_ VGND VPWR VPWR VGND _1018_ _1014_ _1017_ _0976_ sky130_fd_sc_hd__mux2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.i_regbuf\[27\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[27\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[31\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7930_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[21\] clknet_leaf_24_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[21\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7861_ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[16\] clknet_leaf_49_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[16\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6812_ VPWR VGND VGND VPWR _3177_ _3179_ _3175_ _3186_ sky130_fd_sc_hd__o21a_1
X_7792_ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[11\] clknet_leaf_1_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[11\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6743_ VPWR VGND _3123_ _3026_ VPWR VGND sky130_fd_sc_hd__buf_2
X_3955_ VPWR VGND VPWR VGND _0804_ _0807_ _0806_ i_tinyqv.cpu.i_core.i_registers.reg_access\[14\]\[2\]
+ _0668_ _0805_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_42_61 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6674_ VGND VPWR VGND VPWR _3061_ _3057_ _3060_ _3051_ _3029_ sky130_fd_sc_hd__a211o_1
XFILLER_0_9_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5625_ VGND VPWR _0157_ _2301_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_3886_ VPWR VGND VPWR VGND _0637_ i_tinyqv.cpu.i_core.i_registers.reg_access\[5\]\[0\]
+ net58 _0738_ i_tinyqv.cpu.i_core.i_registers.reg_access\[11\]\[0\] sky130_fd_sc_hd__a22o_1
X_8413_ i_tinyqv.cpu.is_alu_imm clknet_leaf_6_clk _0511_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5556_ VPWR VGND _2253_ _2251_ i_uart_rx.cycle_counter\[6\] VPWR VGND sky130_fd_sc_hd__and2_1
X_8344_ i_spi.end_txn_reg clknet_leaf_26_clk _0443_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5487_ _2203_ i_uart_tx.cycle_counter\[0\] i_uart_tx.cycle_counter\[2\] net206 _2197_
+ VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
X_8275_ i_tinyqv.mem.qspi_data_buf\[15\] clknet_leaf_17_clk _0374_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_4507_ VGND VPWR VPWR VGND _1346_ _0752_ _1344_ _0916_ _1345_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_13_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4438_ VGND VPWR VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[1\] i_tinyqv.cpu.i_core.i_shift.a\[30\]
+ _1029_ i_tinyqv.cpu.i_core.i_shift.a\[2\] i_tinyqv.cpu.i_core.i_shift.a\[29\] _1103_
+ _1281_ sky130_fd_sc_hd__mux4_1
X_7226_ VPWR VGND VGND VPWR i_tinyqv.cpu.imm\[23\] _3359_ _3516_ sky130_fd_sc_hd__nor2_1
X_7157_ VPWR VGND VGND VPWR _3368_ i_tinyqv.cpu.instr_data\[1\]\[14\] _3366_ i_tinyqv.cpu.instr_data\[0\]\[14\]
+ _3460_ _3459_ sky130_fd_sc_hd__o221a_2
X_4369_ VPWR VGND VGND VPWR i_tinyqv.cpu.instr_data_start\[17\] _0897_ _1212_ sky130_fd_sc_hd__nor2_1
X_6108_ VGND VPWR VPWR VGND _2622_ i_tinyqv.cpu.i_core.i_shift.a\[30\] _2592_ i_tinyqv.cpu.i_core.i_shift.a\[26\]
+ sky130_fd_sc_hd__mux2_1
X_7088_ VPWR VGND VGND VPWR _3398_ _1478_ _3349_ sky130_fd_sc_hd__or2_1
X_6039_ VGND VPWR _0286_ _2585_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xrebuffer50 VGND VPWR net79 net77 VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_607 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XANTENNA_19 i_tinyqv.mem.q_ctrl.addr\[21\] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_6390_ VGND VPWR _2828_ _2806_ _2829_ _2801_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_5410_ VGND VPWR _1427_ _2140_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_613 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5341_ VPWR VGND VPWR VGND _2077_ net108 _2080_ _0094_ sky130_fd_sc_hd__a21oi_1
X_8060_ i_spi.bits_remaining\[2\] clknet_leaf_25_clk _0195_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_112 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.i_regbuf\[28\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[28\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_495 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5272_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[13\] _2024_ _1880_ sky130_fd_sc_hd__nand2_1
X_7011_ VPWR VGND VGND VPWR _3305_ _3314_ _3329_ sky130_fd_sc_hd__nor2_1
X_4223_ VGND VPWR VPWR VGND _1070_ _1069_ _1050_ _1068_ sky130_fd_sc_hd__mux2_1
X_4154_ VPWR VGND VGND VPWR _1001_ _0983_ _0999_ sky130_fd_sc_hd__nor2_4
X_4085_ VGND VPWR VGND VPWR i_tinyqv.cpu.i_core.imm_lo\[11\] i_tinyqv.cpu.i_core.imm_lo\[10\]
+ i_tinyqv.cpu.i_core.imm_lo\[8\] i_tinyqv.cpu.i_core.imm_lo\[9\] _0932_ sky130_fd_sc_hd__and4bb_1
X_7913_ i_tinyqv.cpu.i_core.i_registers.reg_access\[1\]\[0\] clknet_leaf_39_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[4\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7844_ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[31\] clknet_leaf_1_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[31\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7775_ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[26\] clknet_leaf_53_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[26\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.i_regbuf\[31\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[31\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[3\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4987_ VGND VPWR _0015_ _1751_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6726_ VGND VPWR VPWR VGND _3104_ _3108_ _3107_ sky130_fd_sc_hd__xor2_1
XFILLER_0_46_521 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_3938_ VPWR VGND VPWR VGND net62 i_tinyqv.cpu.i_core.i_registers.reg_access\[6\]\[2\]
+ _0639_ _0790_ i_tinyqv.cpu.i_core.i_registers.reg_access\[13\]\[2\] sky130_fd_sc_hd__a22o_1
X_6657_ VGND VPWR _3045_ _3043_ _3044_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_3869_ VPWR VGND VPWR VGND _0708_ _0720_ _0658_ _0721_ sky130_fd_sc_hd__or3_4
X_5608_ VPWR VGND VGND VPWR i_uart_rx.fsm_state\[1\] _2289_ i_uart_rx.fsm_state\[0\]
+ sky130_fd_sc_hd__nand2_1
X_6588_ VGND VPWR _0434_ _2986_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5539_ VPWR VGND _2242_ net17 VPWR VGND sky130_fd_sc_hd__buf_2
X_8327_ i_tinyqv.cpu.instr_data_in\[15\] clknet_leaf_16_clk _0426_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.i_regbuf\[20\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[20\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[24\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_8258_ i_tinyqv.mem.qspi_data_byte_idx\[0\] clknet_leaf_17_clk _0357_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_7209_ VPWR VGND _3504_ _3503_ _3290_ VPWR VGND sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_21_Left_102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_8189_ i_tinyqv.cpu.i_core.i_shift.a\[8\] clknet_leaf_41_clk _0301_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.i_regbuf\[16\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[16\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[20\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_30_Left_111 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_20_421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_32_270 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_instrret.i_regbuf\[15\] i_tinyqv.cpu.i_core.i_instrret.reg_buf\[15\]
+ i_tinyqv.cpu.i_core.i_instrret.register\[19\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5890_ VGND VPWR VPWR VGND _2491_ _2490_ _2399_ i_spi.data\[3\] sky130_fd_sc_hd__mux2_1
X_4910_ VGND VPWR VPWR VGND _1700_ _1638_ _1696_ i_tinyqv.cpu.i_core.i_registers.reg_access\[2\]\[3\]
+ sky130_fd_sc_hd__mux2_1
X_4841_ VGND VPWR VPWR VGND _1661_ i_tinyqv.cpu.debug_rd\[1\] _1659_ i_tinyqv.cpu.i_core.i_registers.reg_access\[11\]\[1\]
+ sky130_fd_sc_hd__mux2_1
X_7560_ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[3\] clknet_leaf_47_clk _0053_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_96 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4772_ VGND VPWR VPWR VGND _1607_ i_tinyqv.cpu.i_core.cycle_count_wide\[6\] _1604_
+ i_tinyqv.cpu.i_core.time_hi\[2\] sky130_fd_sc_hd__mux2_1
X_6511_ VGND VPWR VGND VPWR _2924_ _2925_ _2923_ _1713_ sky130_fd_sc_hd__o21ba_4
X_7491_ VPWR VGND _2878_ _3725_ _3728_ _3730_ _3729_ VPWR VGND sky130_fd_sc_hd__o31ai_1
X_6442_ VGND VPWR VPWR VGND _2873_ _2872_ _2863_ _1706_ sky130_fd_sc_hd__mux2_1
X_6373_ VPWR VGND VGND VPWR _1707_ _2785_ _2813_ sky130_fd_sc_hd__nor2_1
X_8112_ i_tinyqv.cpu.instr_data\[0\]\[12\] clknet_leaf_9_clk _0224_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5324_ VPWR VGND VGND VPWR _2067_ _2068_ _0089_ sky130_fd_sc_hd__nor2_1
X_8043_ i_debug_uart_tx.data_to_send\[5\] clknet_leaf_28_clk _0178_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_498 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5255_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.multiplier.accum\[14\] _2008_ _2007_
+ sky130_fd_sc_hd__nand2_1
X_4206_ VGND VPWR VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[26\] i_tinyqv.cpu.i_core.i_shift.a\[27\]
+ i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt\[0\] i_tinyqv.cpu.i_core.i_shift.a\[5\]
+ i_tinyqv.cpu.i_core.i_shift.a\[4\] _1029_ _1053_ sky130_fd_sc_hd__mux4_1
XFILLER_0_47_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5186_ VGND VPWR VPWR VGND _1940_ _1942_ _1941_ sky130_fd_sc_hd__xor2_1
X_4137_ VPWR VGND VPWR VGND _0984_ i_tinyqv.cpu.data_addr\[2\] sky130_fd_sc_hd__inv_2
X_4068_ VPWR VGND VGND VPWR _0915_ _0897_ _0914_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_454 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_7827_ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[14\] clknet_leaf_4_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[14\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7758_ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[9\] clknet_leaf_47_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[9\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7689_ i_tinyqv.cpu.i_core.i_registers.reg_access\[10\]\[0\] clknet_leaf_1_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[4\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6709_ VGND VPWR _1752_ _3093_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_470 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.i_regbuf\[21\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[21\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[25\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.i_regbuf\[28\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[28\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_207 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.i_regbuf\[17\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[17\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[21\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_605 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_25_557 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.i_regbuf\[20\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[20\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[24\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_613 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_5040_ VGND VPWR _1801_ _1802_ _1800_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_6991_ VPWR VGND VGND VPWR _3312_ _3291_ _3281_ sky130_fd_sc_hd__nand2_2
X_5942_ VGND VPWR VPWR VGND _2527_ _2526_ _2524_ net314 sky130_fd_sc_hd__mux2_1
XFILLER_0_48_627 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_5873_ VGND VPWR VPWR VGND _2481_ i_tinyqv.cpu.instr_data\[0\]\[13\] _2468_ _1717_
+ sky130_fd_sc_hd__mux2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.i_regbuf\[8\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[8\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[12\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7612_ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[23\] clknet_leaf_2_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[23\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4824_ VGND VPWR VPWR VGND _1651_ i_tinyqv.cpu.debug_rd\[2\] _1648_ i_tinyqv.cpu.i_core.i_registers.reg_access\[13\]\[2\]
+ sky130_fd_sc_hd__mux2_1
X_4755_ VGND VPWR _0896_ _1590_ _0881_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_7543_ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[18\] clknet_leaf_46_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[18\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_630 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_50_94 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4686_ VPWR VGND VGND VPWR i_tinyqv.cpu.instr_write_offset\[2\] _1522_ _1519_ sky130_fd_sc_hd__nand2_1
X_7474_ VPWR VGND _3715_ _3707_ i_tinyqv.cpu.instr_data_start\[20\] VPWR VGND sky130_fd_sc_hd__and2_1
X_6425_ VPWR VGND _2859_ _2858_ _2832_ VPWR VGND sky130_fd_sc_hd__and2_1
X_6356_ VPWR VGND VPWR VGND _1706_ _2797_ i_tinyqv.mem.q_ctrl.fsm_state\[1\] _1707_
+ sky130_fd_sc_hd__or3b_2
X_5307_ VPWR VGND VPWR VGND _0855_ _0924_ _1173_ _1026_ _2054_ sky130_fd_sc_hd__or4_2
X_6287_ VGND VPWR VPWR VGND _2753_ _2316_ _1552_ net275 sky130_fd_sc_hd__mux2_1
X_8026_ i_tinyqv.cpu.instr_data\[3\]\[4\] clknet_leaf_10_clk _0161_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5238_ VGND VPWR _1966_ _1963_ _1992_ _1965_ VPWR VGND sky130_fd_sc_hd__o21ai_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.i_regbuf\[6\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[6\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[10\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5169_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[9\] _1925_ _1880_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_705 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_13_505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_4540_ VPWR VGND VPWR VGND _1357_ _0878_ _1378_ _1379_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_10_clk VGND VPWR clknet_3_2__leaf_clk clknet_leaf_10_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_4471_ VPWR VGND _1310_ _1309_ i_tinyqv.cpu.i_core.i_shift.a\[0\] VPWR VGND sky130_fd_sc_hd__and2_1
X_6210_ VPWR VGND VPWR VGND _0868_ _1536_ _0979_ i_tinyqv.mem.qspi_data_byte_idx\[1\]
+ _2691_ sky130_fd_sc_hd__or4_1
X_7190_ VPWR VGND VGND VPWR _1422_ _1432_ _3487_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6141_ VGND VPWR VPWR VGND _2648_ _2647_ _2642_ _0777_ sky130_fd_sc_hd__mux2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.i_regbuf\[10\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[10\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[14\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6072_ VGND VPWR VPWR VGND _2604_ i_tinyqv.cpu.i_core.i_shift.a\[12\] _2593_ i_tinyqv.cpu.i_core.i_shift.a\[8\]
+ sky130_fd_sc_hd__mux2_1
X_5023_ VGND VPWR VPWR VGND _1783_ _0016_ _1785_ sky130_fd_sc_hd__xor2_1
X_6974_ VGND VPWR VGND VPWR _0510_ i_tinyqv.cpu.is_load _3282_ _3296_ _3205_ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_5925_ VGND VPWR VPWR VGND _2515_ i_tinyqv.cpu.i_core.mepc\[6\] _2504_ i_tinyqv.cpu.i_core.i_shift.a\[10\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_5856_ VGND VPWR _0216_ _2472_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_3_Right_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4807_ VPWR VGND VPWR VGND _1640_ i_tinyqv.cpu.i_core.i_registers.rd\[0\] sky130_fd_sc_hd__inv_2
X_8575_ VGND VPWR i_tinyqv.mem.q_ctrl.spi_ram_b_select uio_out[7] VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_5787_ VPWR VGND VGND VPWR i_spi.spi_select _2422_ _2418_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_598 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_8_576 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_16_365 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4738_ VGND VPWR _1573_ _1571_ _1572_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_7526_ VPWR VGND VGND VPWR _3746_ _3753_ _0605_ sky130_fd_sc_hd__nor2_1
X_7457_ VGND VPWR VGND VPWR _3701_ _2878_ _2732_ net161 _3700_ sky130_fd_sc_hd__a211o_1
X_4669_ VPWR VGND VGND VPWR _1505_ i_tinyqv.cpu.instr_data\[2\]\[12\] _1422_ sky130_fd_sc_hd__or2_1
X_6408_ VPWR VGND VGND VPWR _2837_ _2841_ _2844_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_instrret.i_regbuf\[4\] i_tinyqv.cpu.i_core.i_instrret.reg_buf\[4\]
+ i_tinyqv.cpu.i_core.i_instrret.register\[8\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7388_ VPWR VGND VGND VPWR i_tinyqv.cpu.data_addr\[6\] _2682_ _3642_ _3643_ sky130_fd_sc_hd__o21a_1
X_6339_ VGND VPWR _2781_ _1536_ _2181_ _2678_ VPWR VGND sky130_fd_sc_hd__and3_1
X_8009_ i_uart_rx.recieved_data\[2\] clknet_leaf_19_clk _0144_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_390 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_59_clk VGND VPWR clknet_3_0__leaf_clk clknet_leaf_59_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_0_57_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_3971_ VGND VPWR VGND VPWR _0699_ _0823_ _0655_ sky130_fd_sc_hd__or2b_1
X_5710_ VPWR VGND _2361_ _0989_ i_debug_uart_tx.cycle_counter\[0\] i_debug_uart_tx.cycle_counter\[1\]
+ i_debug_uart_tx.cycle_counter\[2\] VGND VPWR sky130_fd_sc_hd__a31o_1
X_6690_ VPWR VGND VGND VPWR _3075_ _2991_ _2517_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_107 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_5_513 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5641_ VGND VPWR VPWR VGND _2313_ i_tinyqv.cpu.instr_data_in\[5\] _2309_ i_tinyqv.cpu.instr_data\[3\]\[5\]
+ sky130_fd_sc_hd__mux2_1
X_5572_ _2238_ _2264_ _2239_ _2262_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_8360_ i_tinyqv.cpu.instr_data_start\[18\] clknet_leaf_36_clk _0459_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_8291_ i_tinyqv.mem.qspi_data_buf\[31\] clknet_leaf_16_clk _0390_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_4523_ VPWR VGND VPWR VGND _1361_ _0971_ _1358_ _1362_ _0973_ sky130_fd_sc_hd__a22o_1
X_7311_ VGND VPWR _0561_ _3582_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_68_Left_149 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold225 net254 i_tinyqv.cpu.i_core.i_registers.reg_access\[9\]\[1\] VPWR VGND VGND
+ VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 net243 i_tinyqv.cpu.alu_op\[3\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold203 net232 i_tinyqv.cpu.i_core.mepc\[8\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7242_ VGND VPWR VGND VPWR _3526_ _3453_ _3510_ _3330_ _3438_ sky130_fd_sc_hd__a211o_1
Xhold236 net265 i_tinyqv.mem.q_ctrl.nibbles_remaining\[1\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 net276 i_tinyqv.mem.qspi_data_buf\[28\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 net287 i_tinyqv.mem.qspi_data_buf\[29\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 net298 i_tinyqv.cpu.data_addr\[10\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4454_ VPWR VGND VPWR VGND _1294_ _1080_ _1296_ _1297_ sky130_fd_sc_hd__a21oi_1
X_4385_ VPWR VGND VGND VPWR _1228_ _1227_ _1226_ sky130_fd_sc_hd__nor2_4
X_7173_ VGND VPWR _3359_ _3474_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_6124_ VGND VPWR VPWR VGND _2635_ _2634_ _2592_ i_tinyqv.cpu.i_core.i_shift.a\[31\]
+ sky130_fd_sc_hd__mux2_1
X_6055_ VGND VPWR _0293_ _2594_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5006_ VGND VPWR _1768_ _1769_ _1767_ VPWR VGND sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_77_Left_158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6957_ VPWR VGND _3280_ _2151_ _2146_ VPWR VGND sky130_fd_sc_hd__and2_1
X_5908_ VGND VPWR _0237_ _2503_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6888_ VGND VPWR _0470_ _3250_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_416 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5839_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_cycles.rstn _2460_ _2307_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_395 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_8558_ i_tinyqv.cpu.i_core.i_cycles.register\[31\] clknet_leaf_51_clk i_tinyqv.cpu.i_core.i_cycles.reg_buf\[31\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7509_ VGND VPWR _3743_ _2073_ _2079_ _3742_ VPWR VGND sky130_fd_sc_hd__and3_1
X_8489_ i_tinyqv.mem.q_ctrl.addr\[15\] clknet_leaf_32_clk _0587_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.i_regbuf\[10\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[10\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[14\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_67_552 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_cycles.i_regbuf\[29\] i_tinyqv.cpu.i_core.i_cycles.reg_buf\[29\]
+ i_tinyqv.cpu.i_core.i_cycles.register\[1\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4170_ VPWR VGND VGND VPWR _1016_ _1017_ _0979_ sky130_fd_sc_hd__nand2_4
X_7860_ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[15\] clknet_leaf_45_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[15\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6811_ VPWR VGND VPWR VGND _3185_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[26\]
+ sky130_fd_sc_hd__inv_2
X_7791_ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[10\] clknet_leaf_56_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[10\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6742_ VGND VPWR VGND VPWR _0452_ i_tinyqv.cpu.instr_data_start\[11\] _3027_ _3122_
+ _3093_ sky130_fd_sc_hd__o211a_1
X_3954_ VPWR VGND VPWR VGND _0675_ i_tinyqv.cpu.i_core.i_registers.reg_access\[8\]\[2\]
+ net25 _0806_ i_tinyqv.cpu.i_core.i_registers.reg_access\[5\]\[2\] sky130_fd_sc_hd__a22o_1
X_6673_ VPWR VGND VGND VPWR _3051_ _3059_ _3060_ sky130_fd_sc_hd__nor2_1
X_3885_ VPWR VGND VPWR VGND net47 i_tinyqv.cpu.i_core.i_registers.reg_access\[15\]\[0\]
+ net84 _0737_ i_tinyqv.cpu.i_core.i_registers.reg_access\[14\]\[0\] sky130_fd_sc_hd__a22o_1
X_5624_ VPWR VGND VGND VPWR _2301_ _2229_ net9 sky130_fd_sc_hd__or2_1
X_8412_ i_tinyqv.cpu.is_load clknet_leaf_7_clk _0510_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_8343_ i_tinyqv.cpu.pc\[2\] clknet_leaf_22_clk _0442_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_14_633 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5555_ VPWR VGND VGND VPWR _2251_ _2252_ _0136_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_655 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_5486_ VGND VPWR VGND VPWR _0117_ _0991_ _2171_ _2200_ _2202_ sky130_fd_sc_hd__o211a_1
X_8274_ i_tinyqv.mem.qspi_data_buf\[14\] clknet_leaf_14_clk _0373_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_4506_ VGND VPWR _0898_ _1345_ _0784_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_4437_ VGND VPWR VPWR VGND _1279_ _1270_ _1046_ _1280_ _1121_ sky130_fd_sc_hd__a31oi_1
X_7225_ VGND VPWR VGND VPWR _3510_ _3315_ _3514_ _3515_ sky130_fd_sc_hd__o21ba_1
X_7156_ VPWR VGND VPWR VGND i_tinyqv.cpu.instr_data\[3\]\[14\] _3369_ _3459_ _3370_
+ i_tinyqv.cpu.instr_data\[2\]\[14\] _3372_ sky130_fd_sc_hd__a221o_1
X_6107_ VGND VPWR _0318_ _2621_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4368_ VGND VPWR VPWR VGND i_tinyqv.cpu.instr_data_start\[21\] _1211_ _0900_ sky130_fd_sc_hd__xor2_1
X_4299_ VGND VPWR VPWR VGND _1146_ _1085_ _1083_ _1082_ sky130_fd_sc_hd__mux2_1
X_7087_ VGND VPWR _0522_ _3397_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6038_ VGND VPWR VPWR VGND _2585_ i_tinyqv.cpu.instr_data\[1\]\[9\] _2463_ _2318_
+ sky130_fd_sc_hd__mux2_1
Xrebuffer51 VGND VPWR net80 _0655_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7989_ i_uart_tx.cycle_counter\[8\] clknet_leaf_31_clk _0124_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_660 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_496 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_63_28 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5340_ VGND VPWR _2077_ _2079_ _2080_ net108 VPWR VGND sky130_fd_sc_hd__o21ai_1
X_5271_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[12\] _2023_ _1813_ sky130_fd_sc_hd__nand2_1
X_4222_ VGND VPWR VPWR VGND _1069_ i_tinyqv.cpu.i_core.i_shift.a\[21\] _1027_ i_tinyqv.cpu.i_core.i_shift.a\[10\]
+ sky130_fd_sc_hd__mux2_1
X_7010_ VPWR VGND _3328_ _3290_ VPWR VGND sky130_fd_sc_hd__buf_2
X_4153_ VPWR VGND VGND VPWR _1000_ _0999_ _0998_ sky130_fd_sc_hd__nor2_4
X_4084_ VPWR VGND VGND VPWR _0926_ _0930_ _0931_ sky130_fd_sc_hd__nor2_1
X_7912_ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[3\] clknet_leaf_48_clk _0061_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7843_ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[30\] clknet_leaf_3_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[30\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4986_ VGND VPWR VPWR VGND _1751_ _1750_ _1742_ i_debug_uart_tx.uart_tx_data\[7\]
+ sky130_fd_sc_hd__mux2_1
X_7774_ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[25\] clknet_leaf_54_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[25\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_703 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_6725_ _3107_ _3105_ _3106_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_3937_ VPWR VGND VPWR VGND _0637_ i_tinyqv.cpu.i_core.i_registers.reg_access\[10\]\[2\]
+ _0646_ _0789_ i_tinyqv.cpu.i_core.i_registers.reg_access\[11\]\[2\] sky130_fd_sc_hd__a22o_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.i_regbuf\[24\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[24\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[28\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6656_ VPWR VGND VGND VPWR _3021_ _3022_ _3019_ _3044_ sky130_fd_sc_hd__o21a_1
XFILLER_0_6_641 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_3868_ VGND VPWR VGND VPWR net21 net23 _0720_ _0698_ sky130_fd_sc_hd__a21oi_2
X_5607_ VPWR VGND VGND VPWR _2281_ _2287_ _2288_ _0152_ sky130_fd_sc_hd__o21a_1
X_6587_ VGND VPWR VPWR VGND _2986_ i_tinyqv.mem.q_ctrl.delay_cycles_cfg\[2\] _1728_
+ net12 sky130_fd_sc_hd__mux2_1
X_3799_ VPWR VGND VPWR VGND _0644_ _0651_ _0650_ i_tinyqv.cpu.i_core.i_registers.reg_access\[9\]\[3\]
+ _0642_ _0647_ sky130_fd_sc_hd__a2111o_1
X_5538_ VPWR VGND VGND VPWR _2240_ _2238_ _2241_ _1228_ sky130_fd_sc_hd__nor3b_1
X_8326_ i_tinyqv.cpu.instr_data_in\[14\] clknet_leaf_13_clk _0425_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_8257_ i_tinyqv.cpu.i_core.multiplier.accum\[15\] clknet_leaf_42_clk _0356_ VPWR
+ VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5469_ VGND VPWR VGND VPWR _0112_ i_debug_uart_tx.uart_tx_data\[4\] _2169_ _2190_
+ _2182_ sky130_fd_sc_hd__o211a_1
X_7208_ VPWR VGND VPWR VGND i_tinyqv.cpu.instr_data\[0\]\[2\] _3487_ _3503_ _3488_
+ i_tinyqv.cpu.instr_data\[1\]\[2\] _3502_ sky130_fd_sc_hd__a221o_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.i_regbuf\[13\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[13\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[17\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_8188_ i_tinyqv.cpu.i_core.i_shift.a\[7\] clknet_leaf_42_clk _0300_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_7139_ VPWR VGND VPWR VGND _3444_ _3314_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_500 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_52_558 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_4840_ VGND VPWR _0034_ _1660_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_405 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6510_ VPWR VGND VGND VPWR _2916_ _1711_ _2813_ i_tinyqv.mem.q_ctrl.spi_clk_out _2924_
+ _1713_ sky130_fd_sc_hd__o221a_1
X_4771_ VPWR VGND VPWR VGND i_tinyqv.cpu.i_core.mie\[19\] _0944_ _1606_ net19 i_tinyqv.cpu.i_core.mepc\[3\]
+ _1605_ sky130_fd_sc_hd__a221o_1
X_7490_ VPWR VGND VPWR VGND _2878_ net177 _2732_ _3729_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_536 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_6441_ VPWR VGND VGND VPWR _2872_ _1540_ _2867_ _2795_ _2846_ _1706_ sky130_fd_sc_hd__o41a_1
X_6372_ VGND VPWR _0392_ _2812_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8111_ i_tinyqv.cpu.instr_data\[0\]\[11\] clknet_leaf_11_clk _0223_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5323_ VPWR VGND VPWR VGND _2057_ net123 _2060_ _2068_ sky130_fd_sc_hd__a21oi_1
X_8042_ i_debug_uart_tx.data_to_send\[4\] clknet_leaf_28_clk _0177_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5254_ VPWR VGND _2007_ _2006_ _2005_ VPWR VGND sky130_fd_sc_hd__and2_1
X_5185_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[10\] _1941_ _1845_ sky130_fd_sc_hd__nand2_1
X_4205_ VGND VPWR VPWR VGND _1052_ _1051_ i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt\[1\]
+ _1049_ sky130_fd_sc_hd__mux2_1
X_4136_ VGND VPWR VPWR VGND _0966_ _0961_ i_tinyqv.cpu.data_addr\[5\] i_tinyqv.cpu.data_addr\[4\]
+ _0983_ sky130_fd_sc_hd__or4_4
X_4067_ VPWR VGND VPWR VGND _0896_ _0881_ i_tinyqv.cpu.instr_data_start\[16\] _0914_
+ sky130_fd_sc_hd__a21oi_1
Xwire20 VGND VPWR net20 _0736_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_19_500 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7826_ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[13\] clknet_leaf_4_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[13\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.i_regbuf\[25\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[25\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[29\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4969_ VPWR VGND _1741_ _1740_ VPWR VGND sky130_fd_sc_hd__buf_2
X_7757_ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[8\] clknet_leaf_1_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[8\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6708_ VPWR VGND VGND VPWR _3037_ _3092_ _3091_ sky130_fd_sc_hd__nand2_1
X_7688_ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[3\] clknet_leaf_54_clk _0037_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6639_ VGND VPWR VGND VPWR _0441_ _0749_ _3027_ _3030_ _2061_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_493 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.i_regbuf\[14\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[14\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[18\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_8309_ i_tinyqv.mem.q_ctrl.spi_data_oe\[0\] clknet_leaf_15_clk _0408_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_19 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.i_regbuf\[9\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[9\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[13\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.i_regbuf\[13\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[13\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[17\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_669 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_cycles.i_regbuf\[11\] i_tinyqv.cpu.i_core.i_cycles.reg_buf\[11\]
+ i_tinyqv.cpu.i_core.i_cycles.register\[15\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6990_ VGND VPWR VGND VPWR _3311_ net249 _3282_ _0511_ sky130_fd_sc_hd__o21ba_1
X_5941_ VGND VPWR VPWR VGND _2526_ i_tinyqv.cpu.i_core.mepc\[11\] _2106_ _1060_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_34_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5872_ VGND VPWR _0224_ _2480_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4823_ VGND VPWR _0043_ _1650_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7611_ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[22\] clknet_leaf_2_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[22\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4754_ VGND VPWR _0617_ _1589_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_7542_ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[17\] clknet_leaf_54_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[17\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_653 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7473_ VPWR VGND VGND VPWR _3714_ i_tinyqv.cpu.instr_data_start\[20\] _3707_ sky130_fd_sc_hd__or2_1
X_4685_ VGND VPWR VGND VPWR _1519_ _1521_ _1520_ sky130_fd_sc_hd__or2b_1
XFILLER_0_43_355 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6424_ VPWR VGND VPWR VGND _2856_ _1713_ _2855_ _2858_ _2857_ sky130_fd_sc_hd__a22o_1
X_6355_ VPWR VGND VPWR VGND _2796_ i_tinyqv.mem.q_ctrl.read_cycles_count\[0\] sky130_fd_sc_hd__inv_2
X_6286_ VGND VPWR _0366_ _2752_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5306_ VGND VPWR _2053_ _0744_ i_tinyqv.cpu.i_core.is_interrupt _2052_ VPWR VGND
+ sky130_fd_sc_hd__and3_1
X_8025_ i_tinyqv.cpu.instr_data\[3\]\[3\] clknet_leaf_13_clk _0160_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5237_ VGND VPWR VPWR VGND _1989_ _1991_ _1990_ sky130_fd_sc_hd__xor2_1
X_5168_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[8\] _1924_ _1813_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_92 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4119_ VPWR VGND VPWR VGND _0963_ _0965_ _0964_ _0962_ _0966_ sky130_fd_sc_hd__or4_2
X_5099_ VGND VPWR _1313_ _1856_ _1858_ _1854_ VPWR VGND sky130_fd_sc_hd__o21ai_1
Xclone3 VPWR VGND net32 _1638_ VPWR VGND sky130_fd_sc_hd__buf_6
XFILLER_0_39_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_7809_ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[28\] clknet_leaf_2_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[28\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_130 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.i_regbuf\[25\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[25\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[29\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_694 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_4_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_20_65 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_4470_ VGND VPWR VGND VPWR _1309_ i_tinyqv.cpu.i_core.cycle\[0\] _0797_ _0793_ sky130_fd_sc_hd__o21a_2
X_6140_ VPWR VGND VPWR VGND _2647_ _0772_ sky130_fd_sc_hd__inv_2
X_6071_ VGND VPWR _0300_ _2603_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5022_ VPWR VGND _1785_ _1583_ _1321_ _1320_ _1784_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_6973_ VGND VPWR VGND VPWR _3296_ _3288_ _3294_ _3284_ _3295_ sky130_fd_sc_hd__a211o_1
X_5924_ VGND VPWR _0242_ _2514_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5855_ VGND VPWR VPWR VGND _2472_ i_tinyqv.cpu.instr_data\[0\]\[4\] _2469_ i_tinyqv.cpu.instr_data_in\[4\]
+ sky130_fd_sc_hd__mux2_1
X_4806_ VGND VPWR _0053_ _1639_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8574_ VGND VPWR i_tinyqv.mem.q_ctrl.spi_ram_a_select uio_out[6] VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_5786_ VPWR VGND VPWR VGND _2421_ net184 sky130_fd_sc_hd__inv_2
X_4737_ VGND VPWR VGND VPWR _1572_ net76 _0797_ i_tinyqv.cpu.i_core.cycle\[0\] i_tinyqv.cpu.i_core.i_shift.a\[1\]
+ sky130_fd_sc_hd__o211a_1
X_7525_ VGND VPWR _3745_ _2049_ _3753_ net217 VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_152 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_7456_ VPWR VGND VPWR VGND _3700_ _2877_ _3699_ _3017_ _3180_ sky130_fd_sc_hd__a211oi_1
X_4668_ VGND VPWR _1449_ _1504_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_163 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6407_ VGND VPWR VGND VPWR _2843_ i_tinyqv.mem.q_ctrl.nibbles_remaining\[0\] _2842_
+ _0396_ sky130_fd_sc_hd__o21ba_1
X_7387_ VPWR VGND VPWR VGND _3641_ _3012_ _2732_ _3642_ sky130_fd_sc_hd__a21oi_1
X_4599_ VGND VPWR VGND VPWR _1433_ _1430_ _1434_ _1435_ _1429_ sky130_fd_sc_hd__a2bb2o_1
X_6338_ VGND VPWR _0390_ _2780_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6269_ VGND VPWR VPWR VGND _0868_ i_tinyqv.mem.q_ctrl.data_ready i_tinyqv.mem.qspi_data_byte_idx\[1\]
+ _2743_ sky130_fd_sc_hd__or3b_1
X_8008_ i_uart_rx.recieved_data\[1\] clknet_leaf_19_clk _0143_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_13_Right_13 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_15_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_3970_ VGND VPWR VGND VPWR _0822_ _0655_ _0699_ sky130_fd_sc_hd__or2b_4
X_5640_ VGND VPWR _0161_ _2312_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5571_ VGND VPWR VGND VPWR _2262_ _2239_ _2263_ _2238_ sky130_fd_sc_hd__nand3_4
XPHY_EDGE_ROW_22_Right_22 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_25_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4522_ VGND VPWR VPWR VGND _1361_ _1360_ _0979_ _1359_ sky130_fd_sc_hd__mux2_1
X_8290_ i_tinyqv.mem.qspi_data_buf\[30\] clknet_leaf_14_clk _0389_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_325 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7310_ VGND VPWR VPWR VGND _3582_ _3581_ _3395_ _0625_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_111 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xhold226 net255 i_debug_uart_tx.data_to_send\[2\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold204 net233 i_debug_uart_tx.data_to_send\[1\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4453_ VPWR VGND VPWR VGND _1295_ _1091_ _1076_ _1296_ sky130_fd_sc_hd__a21o_1
Xhold215 net244 i_tinyqv.cpu.i_core.mepc\[20\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7241_ VGND VPWR _0548_ _3525_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xhold248 net277 i_tinyqv.mem.data_from_read\[17\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold259 net288 i_tinyqv.cpu.data_addr\[19\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 net266 i_tinyqv.cpu.instr_data\[0\]\[14\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4384_ VGND VPWR VGND VPWR i_uart_rx.fsm_state\[1\] i_uart_rx.fsm_state\[3\] i_uart_rx.fsm_state\[2\]
+ _1227_ sky130_fd_sc_hd__nand3b_4
X_7172_ VPWR VGND VGND VPWR net296 _3360_ _3473_ _0531_ sky130_fd_sc_hd__o21a_1
X_6123_ VGND VPWR VGND VPWR _2634_ _2633_ _1395_ _2064_ sky130_fd_sc_hd__a21bo_1
X_6054_ VGND VPWR VPWR VGND _2594_ i_tinyqv.cpu.i_core.i_shift.a\[4\] _2593_ i_tinyqv.cpu.i_core.i_shift.a\[0\]
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_31_Right_31 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5005_ _1768_ _0636_ _0641_ net72 i_tinyqv.cpu.i_core.i_shift.a\[1\] i_tinyqv.cpu.i_core.cycle\[0\]
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__o311a_1
X_6956_ VGND VPWR VGND VPWR _0509_ net180 _1556_ _1604_ _3205_ sky130_fd_sc_hd__o211a_1
X_5907_ VGND VPWR VPWR VGND _2503_ _2500_ _2502_ i_tinyqv.cpu.data_addr\[0\] sky130_fd_sc_hd__mux2_1
X_6887_ VPWR VGND VGND VPWR _3250_ _3246_ _3249_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5838_ VPWR VGND VGND VPWR _2459_ _2066_ i_tinyqv.cpu.instr_data\[1\]\[0\] sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_40_Right_40 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5769_ VPWR VGND VPWR VGND _2408_ i_spi.bits_remaining\[1\] _2406_ _2409_ _2404_
+ sky130_fd_sc_hd__a22o_1
X_8557_ i_tinyqv.cpu.i_core.i_cycles.register\[30\] clknet_leaf_4_clk i_tinyqv.cpu.i_core.i_cycles.reg_buf\[30\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7508_ VPWR VGND VGND VPWR _3742_ i_tinyqv.cpu.i_core.cycle_count\[3\] _2072_ sky130_fd_sc_hd__or2_1
X_8488_ i_tinyqv.mem.q_ctrl.addr\[14\] clknet_leaf_32_clk _0586_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_12_Left_93 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7439_ VPWR VGND VPWR VGND _3684_ _3005_ _3685_ _0586_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_177 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.i_regbuf\[28\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[28\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_214 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_54_269 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_22_111 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_26_42 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_6810_ VGND VPWR VGND VPWR _0458_ i_tinyqv.cpu.instr_data_start\[17\] _3123_ _3184_
+ _3093_ sky130_fd_sc_hd__o211a_1
X_7790_ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[9\] clknet_leaf_56_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[9\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6741_ VPWR VGND VGND VPWR _3122_ _3029_ _3121_ sky130_fd_sc_hd__or2_1
X_3953_ VGND VPWR VPWR VGND _0805_ _0667_ _0666_ i_tinyqv.cpu.i_core.i_registers.reg_access\[10\]\[2\]
+ _0681_ i_tinyqv.cpu.i_core.i_registers.reg_access\[6\]\[2\] sky130_fd_sc_hd__a32o_1
X_6672_ VGND VPWR VPWR VGND _3059_ _3058_ _2987_ _1205_ sky130_fd_sc_hd__mux2_1
X_3884_ VGND VPWR VGND VPWR _0731_ _0735_ _0736_ _0730_ _0734_ sky130_fd_sc_hd__nor4_2
XFILLER_0_45_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5623_ VGND VPWR _0156_ _2300_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8411_ i_tinyqv.cpu.data_ready_latch clknet_leaf_22_clk _0509_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_8342_ i_tinyqv.cpu.pc\[1\] clknet_leaf_22_clk _0441_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_601 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5554_ VGND VPWR _2249_ _2242_ _2252_ net306 VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_0_5_388 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_14_645 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_14_667 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5485_ VPWR VGND VPWR VGND _2197_ i_uart_tx.cycle_counter\[0\] net206 _2202_ sky130_fd_sc_hd__a21o_1
X_8273_ i_tinyqv.mem.qspi_data_buf\[13\] clknet_leaf_14_clk _0372_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_4505_ VPWR VGND VPWR VGND _0617_ _1338_ _1344_ _1339_ _0689_ _1343_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_689 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_1_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_4436_ VGND VPWR VGND VPWR _1143_ _1278_ _1077_ _1272_ _1274_ _1279_ sky130_fd_sc_hd__a311o_1
X_7224_ VPWR VGND VGND VPWR _3289_ _3514_ _3402_ sky130_fd_sc_hd__nand2_1
X_4367_ VPWR VGND VPWR VGND _0617_ _1201_ _1210_ _1203_ _0691_ _1209_ sky130_fd_sc_hd__a221o_1
X_7155_ VGND VPWR _0529_ _3458_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6106_ VGND VPWR VPWR VGND _2621_ i_tinyqv.cpu.i_core.i_shift.a\[29\] _2592_ i_tinyqv.cpu.i_core.i_shift.a\[25\]
+ sky130_fd_sc_hd__mux2_1
X_4298_ VGND VPWR VPWR VGND _1145_ _1081_ _1083_ _1097_ sky130_fd_sc_hd__mux2_1
X_7086_ VGND VPWR VPWR VGND _3397_ _3394_ _3396_ i_tinyqv.cpu.i_core.imm_lo\[2\] sky130_fd_sc_hd__mux2_1
X_6037_ VGND VPWR _0285_ _2584_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xrebuffer30 VGND VPWR net59 net22 VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xrebuffer41 VGND VPWR net70 i_tinyqv.cpu.i_core.i_registers.rs1\[1\] VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xrebuffer52 VGND VPWR net81 _0798_ VPWR VGND sky130_fd_sc_hd__buf_1
X_7988_ i_uart_tx.cycle_counter\[7\] clknet_leaf_31_clk _0123_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_6939_ VGND VPWR VPWR VGND _0496_ _3274_ _3269_ _1619_ _3275_ net113 sky130_fd_sc_hd__a32o_1
XFILLER_0_49_597 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_51_206 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_47_19 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.i_regbuf\[29\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[29\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[1\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_206 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_23_442 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5270_ VPWR VGND VPWR VGND _2022_ i_tinyqv.cpu.i_core.i_shift.a\[15\] sky130_fd_sc_hd__inv_2
X_4221_ VGND VPWR VPWR VGND _1068_ i_tinyqv.cpu.i_core.i_shift.a\[20\] _1028_ i_tinyqv.cpu.i_core.i_shift.a\[11\]
+ sky130_fd_sc_hd__mux2_1
X_4152_ VPWR VGND VPWR VGND _0999_ i_tinyqv.cpu.data_addr\[2\] _0969_ sky130_fd_sc_hd__or2_2
X_4083_ VPWR VGND VPWR VGND i_tinyqv.cpu.i_core.imm_lo\[2\] i_tinyqv.cpu.i_core.imm_lo\[0\]
+ i_tinyqv.cpu.i_core.imm_lo\[1\] i_tinyqv.cpu.i_core.imm_lo\[3\] _0930_ sky130_fd_sc_hd__or4_1
X_7911_ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[2\] clknet_leaf_5_clk _0060_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7842_ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[29\] clknet_leaf_3_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[29\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4985_ VGND VPWR VPWR VGND _1750_ gpio_out_sel\[7\] _1728_ _1544_ sky130_fd_sc_hd__mux2_1
X_7773_ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[24\] clknet_leaf_0_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[24\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6724_ VPWR VGND VGND VPWR i_tinyqv.cpu.instr_data_start\[10\] _3106_ i_tinyqv.cpu.i_core.imm_lo\[10\]
+ sky130_fd_sc_hd__nand2_1
X_3936_ VPWR VGND VPWR VGND _0613_ _0784_ _0787_ _0788_ sky130_fd_sc_hd__a21oi_1
X_6655_ VPWR VGND VGND VPWR _3041_ _3043_ _3042_ sky130_fd_sc_hd__nand2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.i_regbuf\[17\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[17\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[21\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3867_ VGND VPWR VGND VPWR _0716_ _0718_ _0719_ _0715_ _0717_ sky130_fd_sc_hd__nor4_2
XFILLER_0_33_206 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_5606_ VPWR VGND VPWR VGND _2287_ _2281_ _2229_ _2288_ sky130_fd_sc_hd__a21oi_1
X_6586_ VGND VPWR _0433_ _2985_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_3798_ VPWR VGND VPWR VGND _0649_ i_tinyqv.cpu.i_core.i_registers.reg_access\[1\]\[3\]
+ _0648_ _0650_ i_tinyqv.cpu.i_core.i_registers.reg_access\[7\]\[3\] sky130_fd_sc_hd__a22o_1
X_5537_ VGND VPWR VGND VPWR _2240_ _1728_ _2239_ i_uart_rx.fsm_state\[0\] sky130_fd_sc_hd__o21a_2
X_8325_ i_tinyqv.cpu.instr_data_in\[13\] clknet_leaf_14_clk _0424_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_8256_ i_tinyqv.cpu.i_core.multiplier.accum\[14\] clknet_leaf_43_clk _0355_ VPWR
+ VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5468_ VPWR VGND VGND VPWR _2190_ _2179_ _2189_ sky130_fd_sc_hd__or2_1
X_7207_ VGND VPWR VGND VPWR _3502_ i_tinyqv.cpu.instr_data\[2\]\[2\] _1432_ _1457_
+ _3489_ sky130_fd_sc_hd__o211a_1
X_8187_ i_tinyqv.cpu.i_core.i_shift.a\[6\] clknet_leaf_42_clk _0299_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
X_4419_ VGND VPWR VPWR VGND _1262_ _1084_ _1149_ _1098_ sky130_fd_sc_hd__mux2_1
X_5399_ VPWR VGND VGND VPWR _1483_ _2128_ _2129_ sky130_fd_sc_hd__nor2_1
X_7138_ VPWR VGND VPWR VGND _1491_ _3423_ _3443_ _3441_ _3364_ _3442_ sky130_fd_sc_hd__a221o_1
X_7069_ VPWR VGND VPWR VGND _3348_ _1452_ _3284_ _3381_ _2155_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_191 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_52_548 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_16_707 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_4770_ VPWR VGND VGND VPWR _1604_ _0938_ _1605_ sky130_fd_sc_hd__nor2_1
X_6440_ VGND VPWR VGND VPWR _0401_ i_tinyqv.mem.q_ctrl.fsm_state\[1\] _2863_ _2871_
+ _2832_ sky130_fd_sc_hd__o211a_1
X_6371_ VGND VPWR VPWR VGND _2812_ _2809_ _2811_ i_tinyqv.mem.q_ctrl.read_cycles_count\[0\]
+ sky130_fd_sc_hd__mux2_1
X_5322_ VGND VPWR _2066_ _2067_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_8110_ i_tinyqv.cpu.instr_data\[0\]\[10\] clknet_leaf_4_clk _0222_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_8041_ i_debug_uart_tx.data_to_send\[3\] clknet_leaf_28_clk _0176_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5253_ VPWR VGND VGND VPWR _2006_ _2002_ _2004_ sky130_fd_sc_hd__or2_1
X_5184_ VPWR VGND VGND VPWR _1938_ _1940_ _1939_ sky130_fd_sc_hd__nand2_1
X_4204_ VGND VPWR VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[2\] i_tinyqv.cpu.i_core.i_shift.a\[29\]
+ _1036_ i_tinyqv.cpu.i_core.i_shift.a\[3\] i_tinyqv.cpu.i_core.i_shift.a\[28\] _1050_
+ _1051_ sky130_fd_sc_hd__mux4_1
X_4135_ VPWR VGND _0982_ _0971_ _0752_ VPWR VGND sky130_fd_sc_hd__and2_1
X_4066_ VPWR VGND VGND VPWR _0906_ _0724_ _0905_ _0609_ _0913_ _0912_ sky130_fd_sc_hd__o221a_1
X_7825_ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[12\] clknet_leaf_49_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[12\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4968_ VPWR VGND _1740_ _1725_ net14 VPWR VGND sky130_fd_sc_hd__and2_1
X_7756_ i_tinyqv.cpu.i_core.i_registers.reg_access\[8\]\[3\] clknet_leaf_55_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[7\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.i_regbuf\[18\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[18\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[22\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6707_ VPWR VGND VPWR VGND _3083_ _3039_ _3091_ _2995_ _0911_ _3090_ sky130_fd_sc_hd__a221o_1
X_7687_ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[2\] clknet_leaf_57_clk _0036_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_3919_ VGND VPWR VGND VPWR _0770_ _0769_ i_tinyqv.cpu.i_core.i_registers.reg_access\[10\]\[1\]
+ _0666_ _0667_ _0771_ sky130_fd_sc_hd__a311o_1
X_4899_ VGND VPWR _0064_ _1693_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6638_ VGND VPWR VGND VPWR _3030_ _2995_ _2994_ _1415_ _3029_ sky130_fd_sc_hd__a211o_1
X_8308_ i_tinyqv.mem.q_ctrl.spi_clk_out clknet_leaf_15_clk _0407_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_2
X_6569_ VPWR VGND VGND VPWR _2322_ _2952_ _2975_ _2976_ sky130_fd_sc_hd__o21a_1
XFILLER_0_30_710 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_8239_ i_tinyqv.cpu.i_core.mepc\[10\] clknet_leaf_34_clk _0339_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.i_regbuf\[21\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[21\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[25\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_69_Right_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.i_regbuf\[10\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[10\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[14\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.i_regbuf\[9\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[9\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[13\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_78_Right_78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Left_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_18_21 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xi_tinyqv.cpu.i_core.i_instrret.i_regbuf\[20\] i_tinyqv.cpu.i_core.i_instrret.reg_buf\[20\]
+ i_tinyqv.cpu.i_core.i_instrret.register\[24\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5940_ VGND VPWR _0247_ _2525_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5871_ VGND VPWR VPWR VGND _2480_ i_tinyqv.cpu.instr_data\[0\]\[12\] _2468_ _1712_
+ sky130_fd_sc_hd__mux2_1
X_7610_ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[21\] clknet_leaf_52_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[21\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4822_ VGND VPWR VPWR VGND _1650_ i_tinyqv.cpu.debug_rd\[1\] _1648_ i_tinyqv.cpu.i_core.i_registers.reg_access\[13\]\[1\]
+ sky130_fd_sc_hd__mux2_1
X_7541_ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[16\] clknet_leaf_47_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[16\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4753_ VPWR VGND VGND VPWR _1125_ _1588_ _1587_ sky130_fd_sc_hd__nand2_1
X_7472_ VGND VPWR VPWR VGND _3713_ i_tinyqv.mem.q_ctrl.addr\[16\] _3007_ i_tinyqv.mem.q_ctrl.addr\[20\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_397 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_6423_ VGND VPWR _2857_ _2734_ i_tinyqv.cpu.data_addr\[24\] _2841_ VPWR VGND sky130_fd_sc_hd__and3_1
X_4684_ VPWR VGND _1520_ _1518_ i_tinyqv.mem.instr_active i_tinyqv.cpu.instr_fetch_running
+ _1406_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_6354_ VPWR VGND VPWR VGND i_tinyqv.mem.q_ctrl.nibbles_remaining\[1\] i_tinyqv.mem.q_ctrl.nibbles_remaining\[0\]
+ i_tinyqv.mem.q_ctrl.nibbles_remaining\[2\] _2795_ sky130_fd_sc_hd__or3_4
X_6285_ VGND VPWR VPWR VGND _2752_ i_tinyqv.cpu.instr_data_in\[7\] _2744_ _1721_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_94 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5305_ VPWR VGND _2052_ _2050_ i_tinyqv.cpu.i_core.mip\[17\] i_tinyqv.cpu.i_core.mie\[17\]
+ _2051_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_8024_ i_tinyqv.cpu.instr_data\[3\]\[2\] clknet_leaf_13_clk _0159_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5236_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[12\] _1990_ _1845_ sky130_fd_sc_hd__nand2_1
X_5167_ VGND VPWR VPWR VGND _1921_ _0024_ _1923_ sky130_fd_sc_hd__xor2_1
X_4118_ VPWR VGND VPWR VGND i_tinyqv.cpu.data_addr\[16\] i_tinyqv.cpu.data_addr\[18\]
+ i_tinyqv.cpu.data_addr\[19\] i_tinyqv.cpu.data_addr\[17\] _0965_ sky130_fd_sc_hd__or4_1
X_5098_ VPWR VGND VPWR VGND _1313_ _1856_ _1854_ _1857_ sky130_fd_sc_hd__or3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.i_regbuf\[8\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[8\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[12\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4049_ VPWR VGND _0896_ _0895_ i_tinyqv.cpu.instr_data_start\[14\] VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_38_106 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_7808_ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[27\] clknet_leaf_0_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[27\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7739_ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[22\] clknet_leaf_0_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[22\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_364 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_22_529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_30_584 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.i_regbuf\[22\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[22\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[26\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_426 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.i_regbuf\[11\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[11\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[15\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.i_regbuf\[18\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[18\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[22\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_72_429 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_401 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6070_ VGND VPWR VPWR VGND _2603_ i_tinyqv.cpu.i_core.i_shift.a\[11\] _2593_ _1054_
+ sky130_fd_sc_hd__mux2_1
X_5021_ VPWR VGND _1784_ _1582_ _1580_ VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_45_52 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6972_ VPWR VGND VGND VPWR _3295_ _2147_ _2151_ sky130_fd_sc_hd__nand2_2
X_5923_ VGND VPWR VPWR VGND _2514_ _2513_ _2502_ i_tinyqv.cpu.data_addr\[5\] sky130_fd_sc_hd__mux2_1
X_5854_ VGND VPWR _0215_ _2471_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8573_ VGND VPWR i_tinyqv.mem.q_ctrl.spi_clk_out uio_out[3] VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_4805_ VGND VPWR VPWR VGND _1639_ net32 _1190_ i_tinyqv.cpu.i_core.i_registers.reg_access\[15\]\[3\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5785_ VGND VPWR _0198_ _2420_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_589 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7524_ VPWR VGND VGND VPWR _3745_ _3752_ _0604_ sky130_fd_sc_hd__nor2_1
X_4736_ _1571_ _0636_ _0641_ net71 i_tinyqv.cpu.i_core.i_shift.a\[0\] i_tinyqv.cpu.i_core.cycle\[0\]
+ VPWR VGND VGND VPWR sky130_fd_sc_hd__o311a_1
X_7455_ VPWR VGND VGND VPWR _3697_ _3698_ _3239_ _3699_ sky130_fd_sc_hd__o21a_1
X_4667_ VGND VPWR VPWR VGND _1503_ i_tinyqv.cpu.instr_data\[3\]\[12\] _1449_ i_tinyqv.cpu.instr_data\[1\]\[12\]
+ sky130_fd_sc_hd__mux2_1
X_6406_ VPWR VGND _2843_ _2837_ _2802_ i_tinyqv.mem.q_ctrl.nibbles_remaining\[0\]
+ _2305_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_7386_ VPWR VGND VGND VPWR _3640_ _3067_ _3239_ _3639_ _3641_ sky130_fd_sc_hd__o22a_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.i_regbuf\[4\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[4\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[8\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6337_ VGND VPWR VPWR VGND _2780_ _1721_ _2772_ net261 sky130_fd_sc_hd__mux2_1
X_4598_ VPWR VGND VGND VPWR _1406_ _1409_ _1433_ _1434_ sky130_fd_sc_hd__o21a_1
X_6268_ VGND VPWR _0358_ _2742_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8007_ i_uart_rx.recieved_data\[0\] clknet_leaf_27_clk net202 VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_6199_ VGND VPWR VPWR VGND _0349_ _2221_ _1543_ _2682_ _2679_ _1540_ sky130_fd_sc_hd__o2111a_1
X_5219_ VGND VPWR VPWR VGND _1971_ _0026_ _1973_ sky130_fd_sc_hd__xor2_1
XFILLER_0_34_120 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_5570_ VGND VPWR i_uart_rx.fsm_state\[3\] i_uart_rx.fsm_state\[2\] _2262_ i_uart_rx.fsm_state\[1\]
+ VPWR VGND sky130_fd_sc_hd__o21ai_2
X_4521_ VGND VPWR VPWR VGND _1360_ i_tinyqv.cpu.instr_data_in\[14\] _0838_ i_tinyqv.cpu.instr_data_in\[10\]
+ sky130_fd_sc_hd__mux2_1
Xhold205 VPWR VGND VPWR VGND net234 i_debug_uart_tx.uart_tx_data\[6\] sky130_fd_sc_hd__dlymetal6s2s_1
Xhold216 net245 i_tinyqv.mem.data_from_read\[19\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4452_ VGND VPWR VPWR VGND _1295_ _1157_ _1108_ _1139_ sky130_fd_sc_hd__mux2_1
X_7240_ VGND VPWR VPWR VGND _3525_ _3524_ _3396_ i_tinyqv.cpu.imm\[28\] sky130_fd_sc_hd__mux2_1
Xhold249 net278 i_debug_uart_tx.data_to_send\[7\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 net267 i_tinyqv.mem.qspi_data_buf\[26\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 net256 i_tinyqv.mem.qspi_data_buf\[15\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4383_ VPWR VGND VPWR VGND _1226_ i_uart_rx.fsm_state\[0\] sky130_fd_sc_hd__inv_2
X_7171_ VGND VPWR VGND VPWR _3473_ _3468_ _3472_ _3364_ _3438_ sky130_fd_sc_hd__a211o_1
X_6122_ VGND VPWR VPWR VGND _2633_ _2632_ _1124_ _0652_ sky130_fd_sc_hd__mux2_1
X_6053_ VGND VPWR _2592_ _2593_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_5004_ VGND VPWR VGND VPWR _1767_ net76 _0797_ i_tinyqv.cpu.i_core.cycle\[0\] i_tinyqv.cpu.i_core.i_shift.a\[2\]
+ sky130_fd_sc_hd__o211a_1
X_6955_ VGND VPWR VGND VPWR _0508_ net236 _1387_ _3279_ _3205_ sky130_fd_sc_hd__o211a_1
X_5906_ VPWR VGND _2502_ _2501_ VPWR VGND sky130_fd_sc_hd__buf_4
X_6886_ VGND VPWR VPWR VGND _3249_ i_tinyqv.cpu.i_core.mem_op\[1\] _1761_ i_tinyqv.cpu.data_read_n\[1\]
+ sky130_fd_sc_hd__mux2_1
X_5768_ VPWR VGND VGND VPWR _2402_ _2408_ _2407_ sky130_fd_sc_hd__nand2_1
X_8556_ i_tinyqv.cpu.i_core.i_cycles.register\[29\] clknet_leaf_3_clk i_tinyqv.cpu.i_core.i_cycles.reg_buf\[29\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_8487_ i_tinyqv.mem.q_ctrl.addr\[13\] clknet_leaf_32_clk _0585_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_4719_ VPWR VGND VPWR VGND _1555_ _1404_ sky130_fd_sc_hd__inv_2
X_7507_ VPWR VGND VGND VPWR _2072_ _3741_ _0598_ sky130_fd_sc_hd__nor2_1
X_5699_ VGND VPWR VGND VPWR _2354_ _2336_ _2341_ i_debug_uart_tx.data_to_send\[6\]
+ _2353_ sky130_fd_sc_hd__a211o_1
X_7438_ VPWR VGND VPWR VGND _3008_ i_tinyqv.mem.q_ctrl.addr\[10\] _3007_ _3685_ net315
+ sky130_fd_sc_hd__a22o_1
X_7369_ VPWR VGND VPWR VGND i_tinyqv.cpu.instr_write_offset\[3\] _0884_ i_tinyqv.cpu.instr_data_start\[4\]
+ _3626_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_510 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6740_ VGND VPWR VPWR VGND _3121_ _3120_ _3047_ _3113_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_20 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_3952_ _0804_ _0711_ _0611_ _0620_ _0670_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
X_6671_ VPWR VGND VPWR VGND _3058_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[13\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_18_429 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_3883_ VPWR VGND VPWR VGND net55 i_tinyqv.cpu.i_core.i_registers.reg_access\[6\]\[0\]
+ _0639_ _0735_ i_tinyqv.cpu.i_core.i_registers.reg_access\[7\]\[0\] sky130_fd_sc_hd__a22o_1
X_5622_ VPWR VGND VGND VPWR _2300_ _2229_ net193 sky130_fd_sc_hd__or2_1
X_8410_ i_tinyqv.cpu.data_ready_core clknet_leaf_7_clk _0508_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_5553_ VGND VPWR _2251_ net148 i_uart_rx.cycle_counter\[5\] _2246_ VPWR VGND sky130_fd_sc_hd__and3_1
X_8341_ i_tinyqv.mem.q_ctrl.addr\[3\] clknet_leaf_29_clk _0440_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_4504_ VPWR VGND VGND VPWR _0609_ _1340_ _1342_ _0909_ _1343_ sky130_fd_sc_hd__o22ai_1
X_5484_ VPWR VGND VGND VPWR i_uart_tx.cycle_counter\[0\] _2197_ _2201_ _0116_ sky130_fd_sc_hd__o21a_1
X_8272_ i_tinyqv.mem.qspi_data_buf\[12\] clknet_leaf_14_clk _0371_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_4435_ VPWR VGND VPWR VGND _1275_ _1080_ _1277_ _1278_ sky130_fd_sc_hd__a21oi_1
X_7223_ VPWR VGND VGND VPWR i_tinyqv.cpu.imm\[22\] _3360_ _3513_ _0542_ sky130_fd_sc_hd__o21a_1
X_4366_ VPWR VGND VPWR VGND _0748_ _1205_ _1209_ _1208_ _0689_ _0688_ sky130_fd_sc_hd__a221o_1
X_7154_ VGND VPWR VPWR VGND _3458_ _3457_ _3396_ i_tinyqv.cpu.i_core.imm_lo\[9\] sky130_fd_sc_hd__mux2_1
XFILLER_0_1_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_6105_ VGND VPWR _0317_ _2620_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7085_ VGND VPWR _3395_ _3396_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_4297_ VGND VPWR VGND VPWR _1143_ _1142_ _1077_ _1129_ _1133_ _1144_ sky130_fd_sc_hd__a311o_1
X_6036_ VGND VPWR VPWR VGND _2584_ i_tinyqv.cpu.instr_data\[1\]\[8\] _2463_ _2316_
+ sky130_fd_sc_hd__mux2_1
Xrebuffer20 VGND VPWR net49 _0687_ VPWR VGND sky130_fd_sc_hd__buf_1
Xrebuffer42 VGND VPWR net71 net323 VPWR VGND sky130_fd_sc_hd__buf_1
Xrebuffer53 VGND VPWR net82 _1583_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7987_ i_uart_tx.cycle_counter\[6\] clknet_leaf_31_clk _0122_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_532 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6938_ VGND VPWR VPWR VGND _0495_ _3274_ _3268_ _1619_ _3275_ net115 sky130_fd_sc_hd__a32o_1
XFILLER_0_76_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6869_ VGND VPWR VGND VPWR _3238_ _3039_ _3236_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[31\]
+ _3237_ sky130_fd_sc_hd__a211o_1
XFILLER_0_36_248 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_8539_ i_tinyqv.cpu.i_core.i_cycles.register\[12\] clknet_leaf_51_clk i_tinyqv.cpu.i_core.i_cycles.reg_buf\[12\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_42_218 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_11_605 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_11_638 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_627 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_4220_ VGND VPWR VPWR VGND _1067_ _1066_ i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt\[1\]
+ _1063_ sky130_fd_sc_hd__mux2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.i_regbuf\[25\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[25\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[29\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4151_ VPWR VGND VPWR VGND _0998_ i_tinyqv.cpu.data_addr\[4\] _0967_ sky130_fd_sc_hd__or2_2
X_4082_ VPWR VGND VGND VPWR _0928_ _0926_ _0929_ sky130_fd_sc_hd__nor2_1
X_7910_ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[1\] clknet_leaf_5_clk _0059_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7841_ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[28\] clknet_leaf_48_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[28\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4984_ VPWR VGND VPWR VGND _1741_ net234 _1749_ _0014_ sky130_fd_sc_hd__a21o_1
X_7772_ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[23\] clknet_leaf_58_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[23\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6723_ VPWR VGND VGND VPWR i_tinyqv.cpu.instr_data_start\[10\] i_tinyqv.cpu.i_core.imm_lo\[10\]
+ _3105_ sky130_fd_sc_hd__nor2_1
X_3935_ VPWR VGND VPWR VGND _0786_ i_tinyqv.cpu.instr_data_start\[22\] _0610_ _0787_
+ _0752_ sky130_fd_sc_hd__a22o_1
X_6654_ VPWR VGND VGND VPWR _3042_ i_tinyqv.cpu.instr_data_start\[4\] i_tinyqv.cpu.i_core.imm_lo\[4\]
+ sky130_fd_sc_hd__or2_1
X_5605_ VGND VPWR VPWR VGND _2287_ _2286_ _2284_ _2283_ _1227_ i_uart_rx.fsm_state\[0\]
+ sky130_fd_sc_hd__a32o_1
X_3866_ VPWR VGND VPWR VGND _0681_ i_tinyqv.cpu.i_core.i_registers.reg_access\[5\]\[0\]
+ _0675_ _0718_ i_tinyqv.cpu.i_core.i_registers.reg_access\[6\]\[0\] sky130_fd_sc_hd__a22o_1
X_6585_ VGND VPWR VPWR VGND _2985_ i_tinyqv.mem.q_ctrl.delay_cycles_cfg\[1\] _1728_
+ net11 sky130_fd_sc_hd__mux2_1
X_3797_ VGND VPWR _0624_ _0626_ _0649_ _0627_ _0625_ VPWR VGND sky130_fd_sc_hd__and4b_1
X_5536_ VPWR VGND VPWR VGND i_uart_rx.fsm_state\[2\] i_uart_rx.fsm_state\[1\] i_uart_rx.fsm_state\[3\]
+ _2239_ sky130_fd_sc_hd__or3_4
X_8324_ i_tinyqv.cpu.instr_data_in\[12\] clknet_leaf_13_clk _0423_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5467_ VGND VPWR VPWR VGND _2189_ i_uart_tx.data_to_send\[5\] _2177_ i_uart_tx.data_to_send\[4\]
+ sky130_fd_sc_hd__mux2_1
X_8255_ i_tinyqv.cpu.i_core.multiplier.accum\[13\] clknet_leaf_43_clk _0354_ VPWR
+ VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7206_ VPWR VGND VGND VPWR i_tinyqv.cpu.imm\[17\] _3360_ _3501_ _0537_ sky130_fd_sc_hd__o21a_1
X_4418_ VPWR VGND VGND VPWR _0846_ _1260_ _1261_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_660 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_8186_ i_tinyqv.cpu.i_core.i_shift.a\[5\] clknet_leaf_42_clk _0298_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
X_5398_ VPWR VGND VPWR VGND _2128_ _1426_ _2127_ sky130_fd_sc_hd__or2_2
X_4349_ VGND VPWR VPWR VGND _1193_ debug_rd_r\[3\] debug_register_data i_spi.spi_clk_out
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7137_ VPWR VGND VGND VPWR _3351_ _3398_ _1501_ _3442_ sky130_fd_sc_hd__o21a_1
X_7068_ VPWR VGND VGND VPWR net221 _3360_ _3380_ _0520_ sky130_fd_sc_hd__o21a_1
X_6019_ VGND VPWR _0276_ _2575_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_524 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_9_492 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_9_481 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_cycles.i_regbuf\[8\] i_tinyqv.cpu.i_core.i_cycles.reg_buf\[8\]
+ i_tinyqv.cpu.i_core.i_cycles.register\[12\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_58_19 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_40_clk VGND VPWR clknet_3_5__leaf_clk clknet_leaf_40_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_6370_ VPWR VGND VGND VPWR _2305_ _2811_ _2810_ sky130_fd_sc_hd__nor2_2
XFILLER_0_3_624 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_101 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5321_ VPWR VGND _2066_ _1400_ VPWR VGND sky130_fd_sc_hd__buf_4
X_8040_ i_debug_uart_tx.data_to_send\[2\] clknet_leaf_29_clk _0175_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.i_regbuf\[26\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[26\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[30\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_11_468 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5252_ VPWR VGND VGND VPWR _2002_ _2005_ _2004_ sky130_fd_sc_hd__nand2_1
X_5183_ VPWR VGND VGND VPWR _1907_ _1910_ _1939_ _1937_ sky130_fd_sc_hd__nand3_1
X_4203_ VGND VPWR i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt\[0\] _1050_ VPWR
+ VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_48_63 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4134_ VPWR VGND VPWR VGND _0973_ _0958_ _0971_ _0981_ _0980_ sky130_fd_sc_hd__a22o_1
X_4065_ VPWR VGND VGND VPWR _0912_ _0909_ _0911_ sky130_fd_sc_hd__or2_1
Xwire22 VPWR VGND net22 _0719_ VPWR VGND sky130_fd_sc_hd__buf_2
X_7824_ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[11\] clknet_leaf_52_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[11\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4967_ VPWR VGND VPWR VGND _1727_ i_debug_uart_tx.uart_tx_data\[7\] _1739_ _0007_
+ sky130_fd_sc_hd__a21o_1
X_7755_ i_tinyqv.cpu.i_core.i_registers.reg_access\[8\]\[2\] clknet_leaf_47_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[6\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_31_clk VGND VPWR clknet_3_7__leaf_clk clknet_leaf_31_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_6706_ _3090_ _3089_ net40 VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_7686_ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[1\] clknet_leaf_56_clk _0035_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_3918_ VPWR VGND VPWR VGND _0684_ i_tinyqv.cpu.i_core.i_registers.reg_access\[5\]\[1\]
+ _0675_ _0770_ i_tinyqv.cpu.i_core.i_registers.reg_access\[13\]\[1\] sky130_fd_sc_hd__a22o_1
X_4898_ VGND VPWR VPWR VGND _1693_ _1380_ _1690_ i_tinyqv.cpu.i_core.i_registers.reg_access\[5\]\[2\]
+ sky130_fd_sc_hd__mux2_1
X_3849_ VPWR VGND VGND VPWR _0701_ net80 _0700_ sky130_fd_sc_hd__or2_1
X_6637_ VGND VPWR _3028_ _3029_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_6568_ VGND VPWR VGND VPWR _2975_ _2972_ _2974_ _2914_ _2956_ sky130_fd_sc_hd__a211o_1
X_8307_ i_tinyqv.mem.q_ctrl.spi_flash_select clknet_leaf_16_clk _0406_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5519_ VGND VPWR VPWR VGND _0127_ _2225_ _2224_ _2221_ _2200_ net270 sky130_fd_sc_hd__a32o_1
X_6499_ VGND VPWR VPWR VGND _2913_ i_tinyqv.cpu.data_out\[16\] _2912_ i_tinyqv.cpu.data_out\[24\]
+ sky130_fd_sc_hd__mux2_1
X_8238_ i_tinyqv.cpu.i_core.mepc\[9\] clknet_leaf_40_clk _0338_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_8169_ i_tinyqv.cpu.instr_data\[1\]\[4\] clknet_leaf_10_clk _0281_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.i_regbuf\[14\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[14\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[18\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_611 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_22_clk VGND VPWR clknet_3_3__leaf_clk clknet_leaf_22_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_379 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_instrret.i_regbuf\[13\] i_tinyqv.cpu.i_core.i_instrret.reg_buf\[13\]
+ i_tinyqv.cpu.i_core.i_instrret.register\[17\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5870_ VGND VPWR _0223_ _2479_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4821_ VGND VPWR _0042_ _1649_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_13_clk VGND VPWR clknet_3_2__leaf_clk clknet_leaf_13_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_7540_ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[15\] clknet_leaf_46_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[15\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4752_ VGND VPWR VPWR VGND _1587_ _1163_ _1030_ _1122_ sky130_fd_sc_hd__mux2_1
X_7471_ VGND VPWR VGND VPWR _2733_ _3710_ _3711_ _0591_ _3712_ sky130_fd_sc_hd__a2bb2o_1
X_4683_ _1519_ i_tinyqv.cpu.instr_write_offset\[1\] i_tinyqv.cpu.instr_fetch_running
+ i_tinyqv.mem.instr_active _1518_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
X_6422_ VGND VPWR VGND VPWR _2856_ i_tinyqv.cpu.data_read_n\[0\] _0957_ i_tinyqv.cpu.data_read_n\[1\]
+ _1541_ sky130_fd_sc_hd__a211o_1
XFILLER_0_24_560 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_6353_ VGND VPWR VPWR VGND _2793_ _2791_ _2302_ _2794_ sky130_fd_sc_hd__mux2_2
X_6284_ VGND VPWR _0365_ _2751_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5304_ VGND VPWR _2051_ _0991_ i_tinyqv.cpu.i_core.mie\[19\] _1402_ VPWR VGND sky130_fd_sc_hd__and3_1
X_8023_ i_tinyqv.mem.q_ctrl.stop_txn_reg clknet_leaf_16_clk _0158_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5235_ VPWR VGND VGND VPWR _1987_ _1989_ _1988_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_72 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5166_ VPWR VGND VGND VPWR _1897_ _1923_ _1922_ sky130_fd_sc_hd__nand2_1
X_4117_ VPWR VGND VPWR VGND i_tinyqv.cpu.data_addr\[20\] i_tinyqv.cpu.data_addr\[22\]
+ i_tinyqv.cpu.data_addr\[23\] i_tinyqv.cpu.data_addr\[21\] _0964_ sky130_fd_sc_hd__or4_1
X_5097_ VGND VPWR _1855_ _1856_ _1831_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_4048_ VGND VPWR _0895_ _0726_ i_tinyqv.cpu.instr_data_start\[13\] _0894_ VPWR VGND
+ sky130_fd_sc_hd__and3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.i_regbuf\[30\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[30\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[2\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5999_ VGND VPWR _0266_ _2565_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7807_ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[26\] clknet_leaf_57_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[26\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7738_ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[21\] clknet_leaf_55_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[21\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7669_ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[16\] clknet_leaf_59_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[16\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.i_regbuf\[26\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[26\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[30\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_541 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_30_563 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.i_regbuf\[15\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[15\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[19\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_438 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_53_611 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_29_21 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5020_ VPWR VGND _1783_ _1782_ _1780_ VPWR VGND sky130_fd_sc_hd__xor2_2
Xclkbuf_leaf_2_clk VGND VPWR clknet_3_0__leaf_clk clknet_leaf_2_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_6971_ VPWR VGND VPWR VGND _2135_ _3291_ _3293_ _3294_ sky130_fd_sc_hd__a21o_1
X_5922_ VGND VPWR VPWR VGND _2107_ i_tinyqv.cpu.i_core.mepc\[5\] i_tinyqv.cpu.i_core.i_shift.a\[9\]
+ _2513_ sky130_fd_sc_hd__mux2_2
X_5853_ VGND VPWR VPWR VGND _2471_ net291 _2469_ i_tinyqv.cpu.instr_data_in\[3\] sky130_fd_sc_hd__mux2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.i_regbuf\[6\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[6\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[10\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_641 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_8572_ VGND VPWR i_tinyqv.mem.q_ctrl.spi_flash_select uio_out[0] VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_5784_ VGND VPWR VPWR VGND _2420_ net282 _2415_ i_spi.dc_in sky130_fd_sc_hd__mux2_1
X_4804_ VPWR VGND i_tinyqv.cpu.debug_rd\[3\] _1638_ VPWR VGND sky130_fd_sc_hd__buf_6
X_4735_ VPWR VGND _1570_ _1316_ i_tinyqv.cpu.i_core.multiplier.accum\[2\] VPWR VGND
+ sky130_fd_sc_hd__and2_1
X_7523_ VGND VPWR _3750_ _2049_ _3752_ net176 VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7454_ VPWR VGND VGND VPWR i_tinyqv.cpu.instr_data_start\[17\] _3690_ _3698_ sky130_fd_sc_hd__nor2_1
X_4666_ VPWR VGND VGND VPWR _1502_ _1498_ _1501_ sky130_fd_sc_hd__or2_1
X_6405_ VPWR VGND VGND VPWR _2842_ _2837_ _2841_ sky130_fd_sc_hd__or2_1
X_7385_ VPWR VGND VPWR VGND _3634_ _0883_ i_tinyqv.cpu.was_early_branch _3640_ sky130_fd_sc_hd__a21o_1
X_4597_ VPWR VGND VGND VPWR _1433_ i_tinyqv.cpu.instr_write_offset\[2\] _1422_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_251 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_24_390 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6336_ VGND VPWR _0389_ _2779_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6267_ VGND VPWR _2742_ _2733_ _2181_ _2741_ VPWR VGND sky130_fd_sc_hd__and3_1
X_8006_ i_uart_rx.cycle_counter\[10\] clknet_leaf_30_clk _0141_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_6198_ VPWR VGND _2682_ _2681_ VPWR VGND sky130_fd_sc_hd__buf_4
X_5218_ VPWR VGND VGND VPWR _1945_ _1973_ _1972_ sky130_fd_sc_hd__nand2_1
X_5149_ VGND VPWR _1883_ _1879_ _1906_ _1882_ VPWR VGND sky130_fd_sc_hd__o21ai_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.i_regbuf\[4\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[4\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[8\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_132 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_15_12 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.i_regbuf\[30\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[30\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[2\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_28_Left_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_72_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4520_ VGND VPWR VPWR VGND _1359_ i_tinyqv.mem.qspi_data_buf\[30\] _0974_ i_tinyqv.mem.qspi_data_buf\[26\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_305 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_31_99 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4451_ VGND VPWR VPWR VGND _1294_ _1154_ _1088_ _1158_ sky130_fd_sc_hd__mux2_1
Xhold206 net235 i_tinyqv.cpu.i_core.cycle_count\[3\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold217 net246 i_tinyqv.cpu.i_core.time_hi\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold239 net268 i_tinyqv.cpu.i_core.i_registers.reg_access\[1\]\[1\] VPWR VGND VGND
+ VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7170_ VPWR VGND VGND VPWR _3472_ _3455_ _3471_ sky130_fd_sc_hd__or2_1
Xhold228 net257 i_tinyqv.cpu.imm\[13\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4382_ VPWR VGND VPWR VGND _1225_ _0985_ sky130_fd_sc_hd__inv_2
X_6121_ VGND VPWR VPWR VGND _2632_ _2631_ _2625_ _1569_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_7_Right_7 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6052_ VGND VPWR VGND VPWR _1563_ _1124_ _1031_ _2592_ sky130_fd_sc_hd__a21o_2
XPHY_EDGE_ROW_37_Left_118 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5003_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.multiplier.accum\[3\] _1766_ _1576_
+ sky130_fd_sc_hd__nand2_1
X_6954_ VPWR VGND VPWR VGND _1604_ _1556_ i_tinyqv.cpu.data_ready_latch _3279_ sky130_fd_sc_hd__or3_1
X_5905_ VPWR VGND VGND VPWR _2501_ _1758_ _1400_ sky130_fd_sc_hd__nor2_4
X_6885_ VGND VPWR _0469_ _3248_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_46_Left_127 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5836_ VGND VPWR VGND VPWR _0211_ _0990_ _0991_ net116 _2458_ sky130_fd_sc_hd__a211o_1
X_5767_ VPWR VGND VGND VPWR i_spi.bits_remaining\[1\] _2407_ i_spi.bits_remaining\[0\]
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_633 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_8555_ i_tinyqv.cpu.i_core.i_cycles.register\[28\] clknet_leaf_6_clk i_tinyqv.cpu.i_core.i_cycles.reg_buf\[28\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5698_ VPWR VGND _2353_ _2337_ i_debug_uart_tx.data_to_send\[7\] VPWR VGND sky130_fd_sc_hd__and2_1
X_8486_ i_tinyqv.mem.q_ctrl.addr\[12\] clknet_leaf_33_clk _0584_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_4718_ VGND VPWR VGND VPWR _1553_ _1551_ net6 _1442_ _1410_ net5 _1554_ sky130_fd_sc_hd__mux4_1
X_7506_ VGND VPWR _3739_ _2049_ _3741_ i_tinyqv.cpu.i_core.cycle_count\[2\] VPWR VGND
+ sky130_fd_sc_hd__o21ai_1
X_7437_ VGND VPWR VPWR VGND _3684_ _3683_ _3012_ net111 sky130_fd_sc_hd__mux2_1
X_4649_ VGND VPWR VPWR VGND _1485_ i_tinyqv.cpu.instr_data\[2\]\[15\] net34 i_tinyqv.cpu.instr_data\[0\]\[15\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_636 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.i_regbuf\[29\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[29\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[1\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_146 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7368_ VPWR VGND VGND VPWR _3624_ _3625_ _2732_ sky130_fd_sc_hd__nand2_4
XPHY_EDGE_ROW_55_Left_136 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6319_ VGND VPWR VPWR VGND _2770_ _1721_ _2762_ net285 sky130_fd_sc_hd__mux2_1
X_7299_ VPWR VGND VGND VPWR _3573_ _2143_ _3351_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_544 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_64_Left_145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_73_Left_154 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_31_691 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_26_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_9_107 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_3951_ VPWR VGND VPWR VGND i_tinyqv.cpu.i_core.i_registers.reg_access\[11\]\[2\]
+ _0664_ _0803_ _0680_ i_tinyqv.cpu.i_core.i_registers.reg_access\[9\]\[2\] _0802_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_129 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_6670_ VGND VPWR VPWR VGND _3057_ _3056_ _2991_ _2513_ sky130_fd_sc_hd__mux2_1
X_3882_ _0734_ _0732_ i_tinyqv.cpu.counter\[4\] _0690_ _0733_ VGND VPWR VPWR VGND
+ sky130_fd_sc_hd__and4_1
X_5621_ VGND VPWR VGND VPWR _0155_ _2291_ _2297_ _2298_ _2299_ sky130_fd_sc_hd__o211a_1
X_5552_ VPWR VGND VGND VPWR _2249_ _2250_ _0135_ sky130_fd_sc_hd__nor2_1
X_8340_ i_tinyqv.mem.q_ctrl.addr\[2\] clknet_leaf_33_clk _0439_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_400 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_8271_ i_tinyqv.mem.qspi_data_buf\[11\] clknet_leaf_21_clk _0370_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_4503_ VPWR VGND VGND VPWR _1342_ _0893_ _1341_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_14_625 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_5483_ VPWR VGND VPWR VGND _2200_ _2201_ i_uart_tx.cycle_counter\[0\] _2197_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_1_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_4434_ VPWR VGND VPWR VGND _1276_ _1092_ _1077_ _1277_ sky130_fd_sc_hd__a21o_1
X_7222_ VGND VPWR VGND VPWR _3362_ _3510_ _3328_ _3330_ _3390_ _3513_ sky130_fd_sc_hd__a311o_1
X_4365_ VPWR VGND VGND VPWR _1208_ _1206_ _1207_ sky130_fd_sc_hd__nand2_2
XFILLER_0_1_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_7153_ VPWR VGND VPWR VGND _2165_ _3398_ _3457_ _3453_ _3315_ _3456_ sky130_fd_sc_hd__a221o_1
X_6104_ VGND VPWR VPWR VGND _2620_ i_tinyqv.cpu.i_core.i_shift.a\[24\] _2595_ i_tinyqv.cpu.i_core.i_shift.a\[28\]
+ sky130_fd_sc_hd__mux2_1
X_7084_ VPWR VGND _3395_ _3358_ VPWR VGND sky130_fd_sc_hd__buf_4
X_4296_ VPWR VGND VGND VPWR _1043_ _1047_ _1143_ sky130_fd_sc_hd__nor2_1
X_6035_ VGND VPWR _0284_ _2583_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xrebuffer21 VGND VPWR net50 net49 VPWR VGND sky130_fd_sc_hd__buf_1
Xrebuffer10 VGND VPWR net39 net38 VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xrebuffer54 VGND VPWR net83 _0633_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xrebuffer43 VGND VPWR net72 net71 VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xrebuffer32 VGND VPWR net61 _0668_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7986_ i_uart_tx.cycle_counter\[5\] clknet_leaf_31_clk _0121_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_6937_ VGND VPWR VPWR VGND _0494_ _3274_ _3267_ _1619_ _3275_ net112 sky130_fd_sc_hd__a32o_1
XFILLER_0_49_577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6868_ VPWR VGND VGND VPWR _1442_ _1599_ _2306_ _3237_ sky130_fd_sc_hd__o21a_1
X_5819_ VGND VPWR _0206_ _2446_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6799_ VPWR VGND VPWR VGND _3174_ net203 sky130_fd_sc_hd__inv_2
X_8538_ i_tinyqv.cpu.i_core.i_cycles.register\[11\] clknet_leaf_50_clk i_tinyqv.cpu.i_core.i_cycles.reg_buf\[11\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_8469_ i_tinyqv.cpu.instr_len\[1\] clknet_leaf_7_clk _0567_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_639 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_13_691 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_67_363 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_55_514 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.i_regbuf\[29\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[29\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[1\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_cycles.i_regbuf\[27\] i_tinyqv.cpu.i_core.i_cycles.reg_buf\[27\]
+ i_tinyqv.cpu.i_core.i_cycles.register\[31\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4150_ VGND VPWR _0996_ _0997_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.i_regbuf\[18\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[18\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[22\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4081_ VPWR VGND VPWR VGND i_tinyqv.cpu.i_core.imm_lo\[2\] i_tinyqv.cpu.i_core.imm_lo\[0\]
+ i_tinyqv.cpu.i_core.imm_lo\[3\] _0928_ i_tinyqv.cpu.i_core.imm_lo\[1\] sky130_fd_sc_hd__or4b_1
X_7840_ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[27\] clknet_leaf_5_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[27\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4983_ VGND VPWR _1749_ gpio_out_sel\[6\] _1737_ _1742_ VPWR VGND sky130_fd_sc_hd__and3_1
X_7771_ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[22\] clknet_leaf_53_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[22\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6722_ VPWR VGND VGND VPWR _3095_ _3098_ _3096_ _3104_ sky130_fd_sc_hd__o21a_1
X_3934_ VPWR VGND VPWR VGND i_tinyqv.cpu.instr_data_start\[6\] _0619_ _0786_ _0690_
+ i_tinyqv.cpu.instr_data_start\[10\] _0785_ sky130_fd_sc_hd__a221o_1
X_6653_ VPWR VGND VGND VPWR i_tinyqv.cpu.instr_data_start\[4\] _3041_ i_tinyqv.cpu.i_core.imm_lo\[4\]
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_396 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_3865_ VPWR VGND VPWR VGND _0684_ i_tinyqv.cpu.i_core.i_registers.reg_access\[12\]\[0\]
+ _0674_ _0717_ i_tinyqv.cpu.i_core.i_registers.reg_access\[13\]\[0\] sky130_fd_sc_hd__a22o_1
X_5604_ VPWR VGND VGND VPWR i_uart_rx.rxd_reg\[0\] _2277_ _2286_ _2285_ sky130_fd_sc_hd__nand3_1
XFILLER_0_5_121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6584_ VGND VPWR _0432_ _2984_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_677 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_3796_ VPWR VGND VGND VPWR _0625_ net87 _0624_ _0626_ _0648_ sky130_fd_sc_hd__nor4b_4
X_5535_ VGND VPWR VGND VPWR i_uart_rx.cycle_counter\[8\] _2237_ i_uart_rx.cycle_counter\[9\]
+ _2238_ i_uart_rx.cycle_counter\[10\] sky130_fd_sc_hd__and4bb_4
X_8323_ i_tinyqv.cpu.instr_data_in\[11\] clknet_leaf_16_clk _0422_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5466_ VGND VPWR VGND VPWR _0111_ i_debug_uart_tx.uart_tx_data\[3\] _2169_ _2188_
+ _2182_ sky130_fd_sc_hd__o211a_1
X_8254_ i_tinyqv.cpu.i_core.multiplier.accum\[12\] clknet_leaf_43_clk _0353_ VPWR
+ VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_72 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4417_ VGND VPWR _1260_ _1254_ _1253_ _1259_ VPWR VGND sky130_fd_sc_hd__and3_1
X_7205_ VGND VPWR VGND VPWR _3501_ _3497_ _3500_ _3476_ _3438_ sky130_fd_sc_hd__a211o_1
X_8185_ i_tinyqv.cpu.i_core.i_shift.a\[4\] clknet_leaf_42_clk _0297_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
X_5397_ VPWR VGND VGND VPWR _1420_ _2127_ _2118_ sky130_fd_sc_hd__nand2_1
X_4348_ VPWR VGND uo_out[1] _1192_ VPWR VGND sky130_fd_sc_hd__buf_4
X_7136_ VPWR VGND VGND VPWR _3368_ i_tinyqv.cpu.instr_data\[1\]\[12\] _3366_ i_tinyqv.cpu.instr_data\[0\]\[12\]
+ _3441_ _3440_ sky130_fd_sc_hd__o221a_1
X_4279_ VGND VPWR VPWR VGND _1126_ _1068_ _1103_ _1065_ sky130_fd_sc_hd__mux2_1
X_7067_ VPWR VGND VPWR VGND _3377_ _3379_ _3380_ _3362_ _3376_ sky130_fd_sc_hd__or4b_2
X_6018_ VGND VPWR VPWR VGND _2575_ i_tinyqv.cpu.instr_data\[2\]\[13\] _2562_ _1717_
+ sky130_fd_sc_hd__mux2_1
X_7969_ i_tinyqv.cpu.i_core.i_registers.rd\[2\] clknet_leaf_6_clk _0106_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_70_325 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_3_636 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer1 VGND VPWR net30 i_tinyqv.cpu.i_core.i_registers.rs1\[3\] VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5320_ VPWR VGND VGND VPWR _2065_ _2051_ _2062_ net159 _0088_ _1753_ sky130_fd_sc_hd__o221a_1
X_5251_ VGND VPWR _1977_ _2003_ _2004_ _1976_ VPWR VGND sky130_fd_sc_hd__o21ai_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.i_regbuf\[19\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[19\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[23\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4202_ VGND VPWR VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[30\] i_tinyqv.cpu.i_core.i_shift.a\[31\]
+ i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt\[0\] i_tinyqv.cpu.i_core.i_shift.a\[1\]
+ i_tinyqv.cpu.i_core.i_shift.a\[0\] _1029_ _1049_ sky130_fd_sc_hd__mux4_1
X_5182_ VPWR VGND VPWR VGND _1910_ _1907_ _1937_ _1938_ sky130_fd_sc_hd__a21o_1
X_4133_ VGND VPWR VPWR VGND _0980_ _0976_ _0979_ _0975_ sky130_fd_sc_hd__mux2_1
X_4064_ VPWR VGND VGND VPWR _0911_ _0892_ _0910_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_78_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_7823_ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[10\] clknet_leaf_5_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[10\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7754_ i_tinyqv.cpu.i_core.i_registers.reg_access\[8\]\[1\] clknet_leaf_46_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[5\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5837__1 VPWR VGND VPWR VGND net29 clknet_leaf_18_clk sky130_fd_sc_hd__inv_2
X_4966_ VGND VPWR _1739_ gpio_out\[7\] _1737_ _1730_ VPWR VGND sky130_fd_sc_hd__and3_1
X_6705_ VGND VPWR VPWR VGND _3089_ _3088_ _2990_ _2519_ sky130_fd_sc_hd__mux2_1
X_7685_ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[0\] clknet_leaf_57_clk _0034_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.i_regbuf\[22\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[22\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[26\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4897_ VGND VPWR _0063_ _1692_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_3917_ VPWR VGND VPWR VGND net320 i_tinyqv.cpu.i_core.i_registers.reg_access\[7\]\[1\]
+ _0678_ _0769_ i_tinyqv.cpu.i_core.i_registers.reg_access\[1\]\[1\] sky130_fd_sc_hd__a22o_1
X_6636_ VPWR VGND _3028_ _2306_ _1442_ VPWR VGND sky130_fd_sc_hd__and2_1
X_3848_ VGND VPWR _0699_ _0700_ _0658_ VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_388 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6567_ VGND VPWR VGND VPWR _2974_ i_tinyqv.cpu.data_out\[15\] _2912_ _2929_ _2973_
+ sky130_fd_sc_hd__o211a_1
X_3779_ VGND VPWR VGND VPWR i_tinyqv.cpu.i_core.i_registers.rs1\[0\] i_tinyqv.cpu.i_core.i_registers.rs1\[1\]
+ i_tinyqv.cpu.i_core.i_registers.rs1\[2\] i_tinyqv.cpu.i_core.i_registers.rs1\[3\]
+ _0631_ sky130_fd_sc_hd__and4bb_1
X_8306_ i_tinyqv.mem.q_ctrl.spi_ram_a_select clknet_leaf_17_clk _0405_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5518_ VPWR VGND VGND VPWR _2197_ _2225_ _2174_ sky130_fd_sc_hd__nand2_1
X_6498_ VGND VPWR _2911_ _2912_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_5449_ VPWR VGND VPWR VGND _2175_ _2174_ sky130_fd_sc_hd__inv_2
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.i_regbuf\[11\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[11\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[15\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_8237_ i_tinyqv.cpu.i_core.mepc\[8\] clknet_leaf_40_clk _0337_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_8168_ i_tinyqv.cpu.instr_data\[1\]\[3\] clknet_leaf_13_clk _0280_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_7119_ VPWR VGND VPWR VGND i_tinyqv.cpu.instr_data\[3\]\[10\] _1504_ _3426_ _1461_
+ i_tinyqv.cpu.instr_data\[2\]\[10\] _3371_ sky130_fd_sc_hd__a221o_1
X_8099_ i_debug_uart_tx.resetn net29 net1 VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_4820_ VGND VPWR VPWR VGND _1649_ i_tinyqv.cpu.debug_rd\[0\] _1648_ i_tinyqv.cpu.i_core.i_registers.reg_access\[13\]\[0\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_21 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_4751_ VGND VPWR VGND VPWR _1586_ _1569_ _1585_ _1563_ _1125_ sky130_fd_sc_hd__a211o_1
X_4682_ VGND VPWR _1518_ i_tinyqv.mem.qspi_data_byte_idx\[0\] _0864_ i_tinyqv.mem.q_ctrl.data_ready
+ VPWR VGND sky130_fd_sc_hd__and3_1
X_7470_ VGND VPWR VPWR VGND _3712_ i_tinyqv.mem.q_ctrl.addr\[19\] _3624_ i_tinyqv.mem.q_ctrl.addr\[15\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_76 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_16_528 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_16_539 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_6421_ VGND VPWR VPWR VGND _2840_ _2855_ i_tinyqv.mem.q_ctrl.last_ram_a_sel _2838_
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_43_369 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_12_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_6352_ VPWR VGND VPWR VGND _1711_ _2792_ _2789_ _2793_ sky130_fd_sc_hd__a21o_1
X_6283_ VGND VPWR VPWR VGND _2751_ i_tinyqv.cpu.instr_data_in\[6\] _2744_ _1720_ sky130_fd_sc_hd__mux2_1
X_5303_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.mie\[16\] _2050_ i_tinyqv.cpu.i_core.mip\[16\]
+ sky130_fd_sc_hd__nand2_1
X_8022_ i_uart_rx.rxd_reg\[1\] clknet_leaf_27_clk _0157_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5234_ VPWR VGND VGND VPWR _1957_ _1960_ _1988_ _1986_ sky130_fd_sc_hd__nand3_1
X_5165_ VGND VPWR VGND VPWR _1922_ _1874_ _1871_ _1899_ sky130_fd_sc_hd__a21bo_1
X_4116_ VPWR VGND VPWR VGND i_tinyqv.cpu.data_addr\[8\] i_tinyqv.cpu.data_addr\[10\]
+ i_tinyqv.cpu.data_addr\[11\] i_tinyqv.cpu.data_addr\[9\] _0963_ sky130_fd_sc_hd__or4_1
X_5096_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[6\] _1855_ _1309_ sky130_fd_sc_hd__nand2_1
X_4047_ VPWR VGND _0894_ _0893_ i_tinyqv.cpu.instr_data_start\[11\] VPWR VGND sky130_fd_sc_hd__and2_1
X_7806_ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[25\] clknet_leaf_1_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[25\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5998_ VGND VPWR VPWR VGND _2565_ i_tinyqv.cpu.instr_data\[2\]\[3\] _2563_ i_tinyqv.cpu.instr_data_in\[3\]
+ sky130_fd_sc_hd__mux2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.i_regbuf\[23\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[23\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[27\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4949_ VGND VPWR _1728_ _1729_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_7737_ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[20\] clknet_leaf_59_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[20\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_100 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7668_ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[15\] clknet_leaf_46_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[15\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6619_ VPWR VGND VPWR VGND _3013_ net93 _3009_ _0438_ _3005_ sky130_fd_sc_hd__a22o_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.i_regbuf\[9\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[9\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[13\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_336 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_15_572 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7599_ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[10\] clknet_leaf_2_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[10\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.i_regbuf\[12\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[12\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[16\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.i_regbuf\[19\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[19\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[23\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.i_regbuf\[7\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[7\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[11\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_686 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_52_166 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.i_regbuf\[11\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[11\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[15\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_79 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6970_ VPWR VGND VPWR VGND _3292_ _1483_ _2132_ _3293_ _2118_ sky130_fd_sc_hd__a22o_1
X_5921_ VGND VPWR _0241_ _2512_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5852_ VGND VPWR _0214_ _2470_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8571_ VGND VPWR net1 uio_oe[7] VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_5783_ VGND VPWR _0197_ _2419_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4803_ VGND VPWR VGND VPWR _1638_ _1637_ _1586_ _1034_ _1588_ sky130_fd_sc_hd__a31o_4
X_7522_ VPWR VGND VGND VPWR _3750_ _3751_ _0603_ sky130_fd_sc_hd__nor2_1
X_4734_ VGND VPWR VGND VPWR _1569_ _1175_ _1564_ _0822_ _1568_ sky130_fd_sc_hd__a211o_1
XFILLER_0_9_21 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_7453_ VPWR VGND _3697_ _3690_ i_tinyqv.cpu.instr_data_start\[17\] VPWR VGND sky130_fd_sc_hd__and2_1
X_4665_ VGND VPWR VPWR VGND _1409_ _1500_ _1499_ _1501_ sky130_fd_sc_hd__mux2_2
X_6404_ VPWR VGND VGND VPWR i_tinyqv.mem.q_ctrl.last_ram_a_sel _2838_ _2840_ _2841_
+ sky130_fd_sc_hd__o21a_1
X_7384_ VPWR VGND VGND VPWR _0883_ _3634_ _3639_ sky130_fd_sc_hd__nor2_1
X_4596_ VPWR VGND _1432_ _1409_ VPWR VGND sky130_fd_sc_hd__buf_4
X_6335_ VGND VPWR VPWR VGND _2779_ _1720_ _2772_ net290 sky130_fd_sc_hd__mux2_1
XFILLER_0_3_274 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_8005_ i_uart_rx.cycle_counter\[9\] clknet_leaf_30_clk _0140_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_6266_ VPWR VGND VPWR VGND _2736_ i_tinyqv.mem.qspi_data_byte_idx\[1\] _2735_ _2741_
+ _2740_ sky130_fd_sc_hd__a22o_1
X_6197_ VPWR VGND _2681_ _2680_ VPWR VGND sky130_fd_sc_hd__buf_4
X_5217_ VGND VPWR VGND VPWR _1972_ _1948_ _1919_ _1947_ sky130_fd_sc_hd__a21bo_1
X_5148_ VGND VPWR VPWR VGND _1903_ _1905_ _1904_ sky130_fd_sc_hd__xor2_1
X_5079_ VPWR VGND VGND VPWR _1839_ _1836_ _1837_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_144 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.i_regbuf\[23\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[23\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[27\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4450_ VPWR VGND VGND VPWR _1092_ _1293_ _1292_ sky130_fd_sc_hd__nand2_1
Xhold207 net236 i_tinyqv.cpu.data_ready_core VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 net247 i_uart_rx.cycle_counter\[9\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4381_ VPWR VGND VPWR VGND i_uart_rx.recieved_data\[1\] _0997_ _1224_ uo_out[1] _1001_
+ _0974_ sky130_fd_sc_hd__a221o_1
Xhold229 net258 i_tinyqv.cpu.i_core.mem_op\[1\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6120_ VPWR VGND VPWR VGND _2631_ net49 sky130_fd_sc_hd__inv_2
X_6051_ VGND VPWR _0292_ _2591_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5002_ VGND VPWR VGND VPWR _1315_ _1765_ _1575_ sky130_fd_sc_hd__or2b_1
X_6953_ VPWR VGND VGND VPWR _0505_ _1589_ _0956_ _2087_ _0507_ sky130_fd_sc_hd__o22a_1
XFILLER_0_72_74 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6884_ VPWR VGND VGND VPWR _3248_ _3246_ _3247_ sky130_fd_sc_hd__or2_1
Xclkbuf_3_5__f_clk VGND VPWR VGND VPWR clknet_0_clk clknet_3_5__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_5904_ VGND VPWR VPWR VGND _2500_ i_tinyqv.cpu.i_core.i_shift.a\[4\] _1393_ i_tinyqv.cpu.i_core.mepc\[0\]
+ sky130_fd_sc_hd__mux2_1
X_5835_ VPWR VGND VGND VPWR _2221_ _2458_ _2170_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_589 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5766_ VPWR VGND VGND VPWR _2394_ _2404_ _2406_ sky130_fd_sc_hd__nor2_1
X_8554_ i_tinyqv.cpu.i_core.i_cycles.register\[27\] clknet_leaf_51_clk i_tinyqv.cpu.i_core.i_cycles.reg_buf\[27\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5697_ VGND VPWR VGND VPWR _0178_ i_debug_uart_tx.uart_tx_data\[5\] _2330_ _2352_
+ _2299_ sky130_fd_sc_hd__o211a_1
X_8485_ i_tinyqv.mem.q_ctrl.addr\[11\] clknet_leaf_32_clk _0583_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_4717_ VPWR VGND VGND VPWR i_tinyqv.mem.instr_active _1553_ _1552_ sky130_fd_sc_hd__nand2_1
X_7505_ VPWR VGND VGND VPWR _3739_ _3740_ _0597_ sky130_fd_sc_hd__nor2_1
X_4648_ VGND VPWR VPWR VGND _1484_ i_tinyqv.cpu.instr_data\[3\]\[15\] net35 i_tinyqv.cpu.instr_data\[1\]\[15\]
+ sky130_fd_sc_hd__mux2_1
X_7436_ VPWR VGND VPWR VGND _3680_ _3632_ _3150_ _3683_ _3682_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_7367_ VGND VPWR VGND VPWR net155 _3624_ _1709_ sky130_fd_sc_hd__nand2_8
X_4579_ VPWR VGND VPWR VGND _1415_ _1208_ sky130_fd_sc_hd__inv_2
X_6318_ VGND VPWR _0381_ _2769_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7298_ VGND VPWR VPWR VGND _3570_ _3571_ _3341_ _3572_ sky130_fd_sc_hd__or3_2
X_6249_ _2727_ _1060_ _2694_ _2696_ _2726_ VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_0_50_456 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_10_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold90 net119 i_tinyqv.cpu.data_out\[26\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3950_ VGND VPWR VPWR VGND _0802_ _0670_ _0667_ i_tinyqv.cpu.i_core.i_registers.reg_access\[2\]\[2\]
+ net24 i_tinyqv.cpu.i_core.i_registers.reg_access\[1\]\[2\] sky130_fd_sc_hd__a32o_1
X_3881_ VPWR VGND VGND VPWR _0625_ net324 _0733_ sky130_fd_sc_hd__nor2_1
X_5620_ VPWR VGND _2299_ _1729_ VPWR VGND sky130_fd_sc_hd__buf_2
X_5551_ VGND VPWR _2246_ _2242_ _2250_ net148 VPWR VGND sky130_fd_sc_hd__o21ai_1
X_8270_ i_tinyqv.mem.qspi_data_buf\[10\] clknet_leaf_14_clk _0369_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_4502_ VPWR VGND VPWR VGND _0892_ _0882_ i_tinyqv.cpu.instr_data_start\[10\] _1341_
+ sky130_fd_sc_hd__a21oi_1
X_5482_ VPWR VGND _2200_ _2199_ VPWR VGND sky130_fd_sc_hd__buf_2
X_7221_ VPWR VGND VGND VPWR _3512_ _3474_ i_tinyqv.cpu.imm\[21\] _3510_ _0541_ sky130_fd_sc_hd__o22a_1
XFILLER_0_13_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_4433_ VGND VPWR VPWR VGND _1276_ _1053_ _1088_ _1051_ sky130_fd_sc_hd__mux2_1
X_4364_ VPWR VGND VGND VPWR _1207_ i_tinyqv.cpu.instr_len\[1\] i_tinyqv.cpu.pc\[1\]
+ sky130_fd_sc_hd__or2_1
X_7152_ VGND VPWR VGND VPWR _3456_ _2143_ _3448_ _3299_ _3455_ sky130_fd_sc_hd__a211o_1
XFILLER_0_1_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_4295_ VPWR VGND VPWR VGND _1136_ _1091_ _1141_ _1142_ sky130_fd_sc_hd__a21oi_1
X_6103_ VGND VPWR _0316_ _2619_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7083_ VGND VPWR VGND VPWR _3394_ _2133_ _3388_ _1491_ _3393_ sky130_fd_sc_hd__a211o_1
X_6034_ VGND VPWR VPWR VGND _2583_ i_tinyqv.cpu.instr_data\[1\]\[7\] _2463_ i_tinyqv.cpu.instr_data_in\[7\]
+ sky130_fd_sc_hd__mux2_1
Xrebuffer11 VPWR VGND VPWR VGND net325 _1339_ sky130_fd_sc_hd__dlymetal6s2s_1
X_7985_ i_uart_tx.cycle_counter\[4\] clknet_leaf_32_clk _0120_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_16_Left_97 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xrebuffer55 VGND VPWR net84 _0633_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xrebuffer44 VGND VPWR net73 net71 VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xrebuffer33 VGND VPWR net62 _0628_ VPWR VGND sky130_fd_sc_hd__buf_1
Xrebuffer22 VGND VPWR net51 i_tinyqv.cpu.i_core.i_registers.rs1\[2\] VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_501 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6936_ VGND VPWR VPWR VGND _0493_ _3274_ _3261_ _1619_ _3275_ net129 sky130_fd_sc_hd__a32o_1
XFILLER_0_9_642 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_6867_ VGND VPWR VGND VPWR _3236_ _3040_ _3234_ _3235_ _2993_ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_686 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5818_ _2446_ _2083_ _2445_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_6798_ VGND VPWR VGND VPWR _0457_ i_tinyqv.cpu.instr_data_start\[16\] _3123_ _3173_
+ _3093_ sky130_fd_sc_hd__o211a_1
X_5749_ VGND VPWR VPWR VGND _2391_ net4 _2386_ i_debug_uart_tx.uart_tx_data\[0\] sky130_fd_sc_hd__mux2_1
X_8537_ i_tinyqv.cpu.i_core.cycle_count_wide\[6\] clknet_leaf_5_clk i_tinyqv.cpu.i_core.i_cycles.reg_buf\[10\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_8468_ i_tinyqv.cpu.i_core.i_registers.rs2\[3\] clknet_leaf_52_clk _0566_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_8399_ i_tinyqv.cpu.data_out\[24\] clknet_leaf_20_clk _0497_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_7419_ VPWR VGND VPWR VGND _3632_ _3119_ _3669_ _3666_ _3668_ _2877_ sky130_fd_sc_hd__a221o_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.i_regbuf\[26\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[26\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[30\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_206 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_50_220 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_50_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4080_ VPWR VGND VGND VPWR _0922_ _0926_ _0927_ sky130_fd_sc_hd__nor2_1
X_4982_ VPWR VGND VPWR VGND _1741_ net237 _1748_ _0013_ sky130_fd_sc_hd__a21o_1
X_7770_ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[21\] clknet_leaf_54_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[21\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6721_ VPWR VGND VPWR VGND _3103_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[18\]
+ sky130_fd_sc_hd__inv_2
X_3933_ VPWR VGND VPWR VGND _0617_ net85 _0615_ _0785_ i_tinyqv.cpu.instr_data_start\[14\]
+ sky130_fd_sc_hd__a22o_1
X_6652_ VGND VPWR _1390_ _3040_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_3864_ VPWR VGND VPWR VGND _0680_ i_tinyqv.cpu.i_core.i_registers.reg_access\[14\]\[0\]
+ _0668_ _0716_ i_tinyqv.cpu.i_core.i_registers.reg_access\[9\]\[0\] sky130_fd_sc_hd__a22o_1
X_5603_ VPWR VGND VGND VPWR i_uart_rx.fsm_state\[0\] _1227_ _2285_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_645 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_6583_ VGND VPWR VPWR VGND _2984_ i_tinyqv.mem.q_ctrl.delay_cycles_cfg\[0\] _1737_
+ net10 sky130_fd_sc_hd__mux2_1
X_8322_ i_tinyqv.cpu.instr_data_in\[10\] clknet_leaf_13_clk _0421_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_3795_ VPWR VGND VPWR VGND _0646_ i_tinyqv.cpu.i_core.i_registers.reg_access\[5\]\[3\]
+ _0645_ _0647_ i_tinyqv.cpu.i_core.i_registers.reg_access\[10\]\[3\] sky130_fd_sc_hd__a22o_1
XFILLER_0_42_710 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5534_ VGND VPWR VGND VPWR i_uart_rx.cycle_counter\[7\] i_uart_rx.cycle_counter\[6\]
+ _2235_ _2236_ _2237_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_78_51 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_8253_ i_tinyqv.mem.qspi_write_done clknet_leaf_17_clk _0082_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_5465_ VPWR VGND VGND VPWR _2188_ _2179_ _2187_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_264 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_361 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_8184_ i_tinyqv.cpu.i_core.i_shift.a\[3\] clknet_leaf_41_clk _0296_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
X_4416_ VGND VPWR VPWR VGND _1259_ _1257_ _1258_ _0831_ _1177_ sky130_fd_sc_hd__o2bb2a_1
X_7204_ VPWR VGND VPWR VGND _3465_ _3364_ _3499_ _3500_ sky130_fd_sc_hd__a21o_1
X_5396_ VPWR VGND VGND VPWR _2125_ _2126_ _2122_ sky130_fd_sc_hd__nor2_2
X_7135_ VPWR VGND VPWR VGND i_tinyqv.cpu.instr_data\[3\]\[12\] _3369_ _3440_ _3370_
+ i_tinyqv.cpu.instr_data\[2\]\[12\] _3372_ sky130_fd_sc_hd__a221o_1
X_4347_ VGND VPWR VPWR VGND _1192_ gpio_out\[1\] gpio_out_sel\[1\] i_uart_rx.uart_rts
+ sky130_fd_sc_hd__mux2_1
X_4278_ VPWR VGND VGND VPWR _1031_ _1125_ _1124_ sky130_fd_sc_hd__nor2_2
X_7066_ VPWR VGND VGND VPWR _3346_ _3313_ _3342_ _1490_ _3379_ _3378_ sky130_fd_sc_hd__o221a_1
X_6017_ VGND VPWR _0275_ _2574_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7968_ i_tinyqv.cpu.i_core.i_registers.rd\[1\] clknet_leaf_5_clk _0105_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_6919_ VGND VPWR VPWR VGND _0481_ _3265_ _3261_ _0691_ _3270_ net186 sky130_fd_sc_hd__a32o_1
X_7899_ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[22\] clknet_leaf_3_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[22\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_294 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_20_437 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.i_regbuf\[27\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[27\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[31\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_55_367 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_24_710 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xrebuffer2 VPWR VGND net31 _1546_ VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_0_3_648 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_5250_ VPWR VGND VGND VPWR _2003_ _1951_ _1998_ sky130_fd_sc_hd__or2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.i_regbuf\[30\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[30\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[2\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4201_ VPWR VGND VPWR VGND _1048_ _1043_ _1047_ sky130_fd_sc_hd__or2_2
XFILLER_0_48_21 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5181_ VPWR VGND VGND VPWR _1935_ _1937_ _1936_ sky130_fd_sc_hd__nand2_1
X_4132_ VGND VPWR VPWR VGND _0977_ i_tinyqv.mem.qspi_write_done _0979_ _0978_ sky130_fd_sc_hd__o21a_4
X_4063_ VPWR VGND VGND VPWR i_tinyqv.cpu.instr_data_start\[8\] _0891_ _0910_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_45 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7822_ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[9\] clknet_leaf_5_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[9\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4965_ VPWR VGND VPWR VGND _1727_ net234 _1738_ _0006_ sky130_fd_sc_hd__a21o_1
X_7753_ i_tinyqv.cpu.i_core.i_registers.reg_access\[8\]\[0\] clknet_leaf_57_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[4\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6704_ VGND VPWR _3087_ _3088_ _3086_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_3916_ VPWR VGND VPWR VGND i_tinyqv.cpu.i_core.i_registers.reg_access\[11\]\[1\]
+ _0664_ _0768_ _0681_ i_tinyqv.cpu.i_core.i_registers.reg_access\[6\]\[1\] _0767_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_80_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7684_ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[31\] clknet_leaf_47_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[31\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4896_ VGND VPWR VPWR VGND _1692_ _1303_ _1690_ i_tinyqv.cpu.i_core.i_registers.reg_access\[5\]\[1\]
+ sky130_fd_sc_hd__mux2_1
X_6635_ VGND VPWR _3026_ _3027_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.i_regbuf\[15\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[15\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[19\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_570 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_3847_ VGND VPWR VPWR VGND _0699_ _0698_ _0697_ _0687_ sky130_fd_sc_hd__mux2_4
X_6566_ VPWR VGND VGND VPWR _2973_ i_debug_uart_tx.uart_tx_data\[7\] _2909_ sky130_fd_sc_hd__or2_1
X_3778_ VGND VPWR VGND VPWR i_tinyqv.cpu.counter\[2\] i_tinyqv.cpu.counter\[4\] _0614_
+ _0630_ sky130_fd_sc_hd__nand3b_2
X_8305_ i_tinyqv.mem.q_ctrl.spi_ram_b_select clknet_leaf_16_clk _0404_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5517_ VPWR VGND VPWR VGND _2223_ _0990_ _2179_ _2224_ sky130_fd_sc_hd__a21o_1
X_6497_ VPWR VGND VGND VPWR _2906_ _2911_ _2907_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_297 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_8236_ i_tinyqv.cpu.i_core.mepc\[7\] clknet_leaf_35_clk _0336_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_5448_ VPWR VGND VPWR VGND _2171_ _2173_ _2172_ i_uart_tx.cycle_counter\[2\] _2174_
+ sky130_fd_sc_hd__or4_1
XFILLER_0_2_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_8167_ i_tinyqv.cpu.instr_data\[1\]\[2\] clknet_leaf_13_clk _0279_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5379_ VGND VPWR _0101_ _2111_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8098_ i_tinyqv.cpu.i_core.interrupt_req\[1\] clknet_leaf_18_clk net3 VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_7118_ VPWR VGND VGND VPWR _1507_ _3346_ _3425_ sky130_fd_sc_hd__nor2_1
X_7049_ VPWR VGND _3362_ _3361_ VPWR VGND sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_29_Right_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Right_38 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Right_47 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_56_Right_56 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4750_ VPWR VGND VGND VPWR _1563_ _1584_ _1585_ sky130_fd_sc_hd__nor2_1
X_4681_ VPWR VGND _1517_ net33 _1387_ _1437_ i_tinyqv.cpu.instr_fetch_running VGND
+ VPWR sky130_fd_sc_hd__a31o_1
X_6420_ VGND VPWR VGND VPWR _0398_ i_tinyqv.mem.q_ctrl.nibbles_remaining\[2\] _2842_
+ _2854_ _2832_ sky130_fd_sc_hd__o211a_1
X_6351_ VPWR VGND VPWR VGND _2792_ i_tinyqv.mem.q_ctrl.is_writing sky130_fd_sc_hd__inv_2
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.i_regbuf\[31\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[31\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[3\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5302_ VGND VPWR VPWR VGND _0086_ _2049_ _1755_ _0862_ _1387_ i_tinyqv.cpu.i_core.cycle\[1\]
+ sky130_fd_sc_hd__o2111a_1
X_6282_ VGND VPWR _0364_ _2750_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8021_ i_uart_rx.rxd_reg\[0\] clknet_leaf_27_clk _0156_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_65_Right_65 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5233_ VPWR VGND VPWR VGND _1960_ _1957_ _1986_ _1987_ sky130_fd_sc_hd__a21o_1
X_5164_ VPWR VGND _1921_ _1920_ _1919_ VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_75_52 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4115_ VPWR VGND VPWR VGND i_tinyqv.cpu.data_addr\[12\] i_tinyqv.cpu.data_addr\[14\]
+ i_tinyqv.cpu.data_addr\[15\] i_tinyqv.cpu.data_addr\[13\] _0962_ sky130_fd_sc_hd__or4_1
X_5095_ VPWR VGND VPWR VGND _1854_ i_tinyqv.cpu.i_core.i_shift.a\[8\] sky130_fd_sc_hd__inv_2
X_4046_ VGND VPWR _0893_ _0882_ i_tinyqv.cpu.instr_data_start\[10\] _0892_ VPWR VGND
+ sky130_fd_sc_hd__and3_1
Xclone7 VPWR VGND VGND VPWR _1410_ _1339_ _1411_ net36 sky130_fd_sc_hd__o21a_1
X_7805_ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[24\] clknet_leaf_2_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[24\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_74_Right_74 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5997_ VGND VPWR _0265_ _2564_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4948_ VPWR VGND _1728_ i_debug_uart_tx.resetn VPWR VGND sky130_fd_sc_hd__buf_4
X_7736_ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[19\] clknet_leaf_53_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[19\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.i_regbuf\[16\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[16\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[20\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7667_ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[14\] clknet_leaf_58_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[14\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4879_ VGND VPWR _0071_ _1682_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_676 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_6618_ VGND VPWR VPWR VGND _3013_ _3011_ _3012_ i_tinyqv.cpu.data_addr\[1\] sky130_fd_sc_hd__mux2_1
XFILLER_0_46_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7598_ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[9\] clknet_leaf_53_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[9\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6549_ VGND VPWR VPWR VGND _2959_ _1712_ _2925_ _2958_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_595 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_8219_ i_tinyqv.cpu.i_core.multiplier.accum\[2\] clknet_leaf_42_clk _0020_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.i_regbuf\[9\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[9\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[13\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Left_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_37_153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_52_112 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_80_487 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.i_regbuf\[7\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[7\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[11\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5920_ VGND VPWR VPWR VGND _2512_ _2511_ _2502_ i_tinyqv.cpu.data_addr\[4\] sky130_fd_sc_hd__mux2_1
X_5851_ VGND VPWR VPWR VGND _2470_ i_tinyqv.cpu.instr_data\[0\]\[2\] _2469_ i_tinyqv.cpu.instr_data_in\[2\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_8570_ VGND VPWR net1 uio_oe[6] VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_5782_ VGND VPWR _2419_ _2417_ _2181_ _2418_ VPWR VGND sky130_fd_sc_hd__and3_1
X_4802_ VPWR VGND VPWR VGND _1614_ _0878_ _1637_ _1636_ _1025_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_71_410 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7521_ VGND VPWR _3744_ _2049_ _3751_ net92 VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_0_28_175 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4733_ VPWR VGND VGND VPWR _0824_ _1177_ _1567_ _1173_ _1568_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_71_432 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_7452_ VGND VPWR _0588_ _3696_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6403_ VPWR VGND VGND VPWR _2839_ _2840_ _2732_ sky130_fd_sc_hd__nor2_2
X_4664_ VGND VPWR VPWR VGND _1500_ i_tinyqv.cpu.instr_data\[2\]\[9\] _1449_ i_tinyqv.cpu.instr_data\[0\]\[9\]
+ sky130_fd_sc_hd__mux2_1
X_7383_ VPWR VGND VGND VPWR _3638_ _3625_ net305 _3637_ _0577_ sky130_fd_sc_hd__o22a_1
X_4595_ _1431_ _1406_ _1409_ _1427_ _1430_ VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_0_9_88 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6334_ VGND VPWR _0388_ _2778_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6265_ VGND VPWR _0868_ _2739_ _2740_ _0864_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_8004_ i_uart_rx.cycle_counter\[8\] clknet_leaf_30_clk _0139_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_5216_ VPWR VGND _1971_ _1970_ _1969_ VPWR VGND sky130_fd_sc_hd__and2_1
X_6196_ VPWR VGND VGND VPWR _2680_ i_tinyqv.mem.instr_active _2679_ sky130_fd_sc_hd__or2_1
X_5147_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[10\] _1904_ _1167_ sky130_fd_sc_hd__nand2_1
X_5078_ VPWR VGND VGND VPWR _1836_ _1838_ _1837_ sky130_fd_sc_hd__nand2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.i_regbuf\[6\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[6\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[10\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4029_ VGND VPWR _0876_ uo_out[4] VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_7719_ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[2\] clknet_leaf_56_clk _0032_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_186 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.i_regbuf\[31\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[31\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[3\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.i_regbuf\[20\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[20\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[24\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.i_regbuf\[16\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[16\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[20\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_476 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold208 net237 i_debug_uart_tx.uart_tx_data\[5\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4380_ VPWR VGND VPWR VGND _1222_ _0971_ _1219_ _1223_ _0973_ sky130_fd_sc_hd__a22o_1
Xhold219 net248 i_tinyqv.cpu.i_core.i_cycles.cy VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_384 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_6050_ VGND VPWR VPWR VGND _2591_ i_tinyqv.cpu.instr_data\[1\]\[15\] _2462_ _1721_
+ sky130_fd_sc_hd__mux2_1
X_5001_ VPWR VGND VGND VPWR _1753_ _1760_ _1764_ _0028_ sky130_fd_sc_hd__o21a_1
X_6952_ VGND VPWR _0506_ _3278_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5903_ VGND VPWR _0236_ _2499_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6883_ VGND VPWR VPWR VGND _3247_ i_tinyqv.cpu.i_core.mem_op\[0\] _1761_ i_tinyqv.cpu.data_read_n\[0\]
+ sky130_fd_sc_hd__mux2_1
X_5834_ VPWR VGND VGND VPWR _2083_ _2457_ _0210_ sky130_fd_sc_hd__nor2_1
X_5765_ VGND VPWR VGND VPWR _0193_ net239 _2404_ _2405_ _2299_ sky130_fd_sc_hd__o211a_1
X_8553_ i_tinyqv.cpu.i_core.i_cycles.register\[26\] clknet_leaf_4_clk i_tinyqv.cpu.i_core.i_cycles.reg_buf\[26\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5696_ VGND VPWR VGND VPWR _2352_ _2336_ _2341_ i_debug_uart_tx.data_to_send\[5\]
+ _2351_ sky130_fd_sc_hd__a211o_1
X_8484_ i_tinyqv.mem.q_ctrl.addr\[10\] clknet_leaf_32_clk _0582_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_4716_ VPWR VGND _1552_ _1518_ VPWR VGND sky130_fd_sc_hd__buf_4
X_7504_ VGND VPWR _2071_ _2049_ _3740_ net121 VPWR VGND sky130_fd_sc_hd__o21ai_1
X_7435_ VPWR VGND VGND VPWR _3010_ _3681_ _3682_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_90 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_4647_ VPWR VGND _1483_ _1482_ VPWR VGND sky130_fd_sc_hd__buf_4
X_7366_ VGND VPWR _0575_ _3623_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_573 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_6317_ VGND VPWR VPWR VGND _2769_ _1720_ _2762_ i_tinyqv.mem.data_from_read\[22\]
+ sky130_fd_sc_hd__mux2_1
X_4578_ VGND VPWR _1412_ _1414_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_7297_ VPWR VGND VPWR VGND _3337_ _3353_ _2121_ _3571_ sky130_fd_sc_hd__or3_1
X_6248_ VPWR VGND VPWR VGND _2726_ _2719_ sky130_fd_sc_hd__inv_2
X_6179_ VGND VPWR _0341_ _2670_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xhold80 net109 i_tinyqv.cpu.data_out\[29\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 net120 i_tinyqv.cpu.data_out\[30\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3880_ VPWR VGND _0732_ _0624_ _0627_ VPWR VGND sky130_fd_sc_hd__and2_1
X_5550_ VPWR VGND _2249_ _2246_ net148 VPWR VGND sky130_fd_sc_hd__and2_1
X_5481_ VPWR VGND VGND VPWR _2198_ _2175_ _2199_ sky130_fd_sc_hd__nor2_1
X_4501_ VGND VPWR _0890_ _1340_ _0883_ VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_424 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_4432_ VGND VPWR VPWR VGND _1275_ _1104_ _1149_ _1055_ sky130_fd_sc_hd__mux2_1
X_7220_ VPWR VGND _3512_ _3384_ _3330_ _3328_ _3362_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_4363_ VPWR VGND VGND VPWR _1206_ i_tinyqv.cpu.instr_len\[1\] i_tinyqv.cpu.pc\[1\]
+ sky130_fd_sc_hd__nand2_2
X_7151_ VPWR VGND VPWR VGND _3454_ _3309_ _1507_ _3455_ sky130_fd_sc_hd__a21oi_1
X_4294_ VPWR VGND VPWR VGND _1140_ _1080_ _1076_ _1141_ sky130_fd_sc_hd__a21o_1
X_6102_ VGND VPWR VPWR VGND _2619_ i_tinyqv.cpu.i_core.i_shift.a\[23\] _2595_ i_tinyqv.cpu.i_core.i_shift.a\[27\]
+ sky130_fd_sc_hd__mux2_1
X_7082_ VPWR VGND VPWR VGND _1501_ _3350_ _3393_ _3363_ _3391_ _3392_ sky130_fd_sc_hd__a221o_1
X_6033_ VGND VPWR _0283_ _2582_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xrebuffer12 VGND VPWR net41 _0652_ VPWR VGND sky130_fd_sc_hd__buf_1
X_7984_ i_uart_tx.cycle_counter\[3\] clknet_leaf_32_clk _0119_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xrebuffer34 VGND VPWR net63 net62 VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xrebuffer45 VGND VPWR net74 _0631_ VPWR VGND sky130_fd_sc_hd__buf_1
Xrebuffer23 VGND VPWR net52 i_tinyqv.cpu.i_core.i_registers.rs1\[2\] VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6935_ VPWR VGND VGND VPWR _3275_ _2081_ _0854_ sky130_fd_sc_hd__or2_1
Xrebuffer56 VGND VPWR i_tinyqv.cpu.pc\[2\] net85 VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_6866_ VPWR VGND VGND VPWR _3235_ _2991_ _2550_ sky130_fd_sc_hd__or2_1
X_5817_ VPWR VGND VPWR VGND _2445_ _0916_ _2441_ _2442_ i_tinyqv.cpu.i_core.mip\[16\]
+ _2444_ sky130_fd_sc_hd__o32a_1
X_6797_ VPWR VGND VGND VPWR _3037_ _3173_ _3172_ sky130_fd_sc_hd__nand2_1
X_5748_ VGND VPWR _0191_ _2390_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8536_ i_tinyqv.cpu.i_core.cycle_count_wide\[5\] clknet_leaf_6_clk i_tinyqv.cpu.i_core.i_cycles.reg_buf\[9\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_498 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5679_ _2328_ _0969_ _2340_ _2339_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_8467_ i_tinyqv.cpu.i_core.i_registers.rs2\[2\] clknet_leaf_52_clk _0565_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_8398_ i_tinyqv.cpu.data_out\[23\] clknet_leaf_20_clk _0496_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_7418_ VPWR VGND VGND VPWR _3010_ _3667_ _3668_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_468 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7349_ VPWR VGND _3612_ i_tinyqv.cpu.additional_mem_ops\[0\] i_tinyqv.cpu.additional_mem_ops\[1\]
+ VPWR VGND sky130_fd_sc_hd__and2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.i_regbuf\[19\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[19\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[23\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_52_clk VGND VPWR clknet_3_1__leaf_clk clknet_leaf_52_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_0_23_468 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_37_12 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xi_tinyqv.cpu.i_core.i_instrret.i_regbuf\[29\] i_tinyqv.cpu.i_core.i_instrret.reg_buf\[29\]
+ i_tinyqv.cpu.i_core.i_instrret.register\[1\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4981_ VGND VPWR _1748_ gpio_out_sel\[5\] _1737_ _1742_ VPWR VGND sky130_fd_sc_hd__and3_1
X_6720_ VGND VPWR VGND VPWR _0450_ _0882_ _3027_ _3102_ _3093_ sky130_fd_sc_hd__o211a_1
X_3932_ VGND VPWR i_tinyqv.cpu.instr_data_start\[18\] _0784_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_43_clk VGND VPWR clknet_3_5__leaf_clk clknet_leaf_43_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_6651_ VGND VPWR _2987_ _3039_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_3863_ VGND VPWR _0715_ _0666_ i_tinyqv.cpu.i_core.i_registers.reg_access\[10\]\[0\]
+ _0667_ VPWR VGND sky130_fd_sc_hd__and3_1
X_5602_ _2284_ i_uart_rx.fsm_state\[0\] i_uart_rx.rxd_reg\[0\] _2239_ _2280_ VPWR
+ VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_6582_ VGND VPWR _0431_ _2983_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5533_ VPWR VGND _2236_ i_uart_rx.cycle_counter\[1\] net91 VPWR VGND sky130_fd_sc_hd__and2_1
X_8321_ i_tinyqv.cpu.instr_data_in\[9\] clknet_leaf_14_clk _0420_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_3794_ VGND VPWR VGND VPWR i_tinyqv.cpu.i_core.i_registers.rs1\[0\] i_tinyqv.cpu.i_core.i_registers.rs1\[2\]
+ i_tinyqv.cpu.i_core.i_registers.rs1\[3\] i_tinyqv.cpu.i_core.i_registers.rs1\[1\]
+ _0646_ sky130_fd_sc_hd__and4bb_1
X_8252_ i_tinyqv.mem.data_stall clknet_leaf_17_clk _0352_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5464_ VGND VPWR VPWR VGND _2187_ i_uart_tx.data_to_send\[4\] _2177_ i_uart_tx.data_to_send\[3\]
+ sky130_fd_sc_hd__mux2_1
X_8183_ i_tinyqv.cpu.i_core.i_shift.a\[2\] clknet_leaf_41_clk _0295_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
X_4415_ VPWR VGND VPWR VGND _1256_ _1255_ _1173_ _1258_ sky130_fd_sc_hd__a21oi_1
X_5395_ VPWR VGND VGND VPWR _2123_ _2125_ _2124_ sky130_fd_sc_hd__nand2_1
X_7203_ VPWR VGND VGND VPWR _3499_ _3470_ _3498_ sky130_fd_sc_hd__or2_1
X_7134_ VPWR VGND VGND VPWR net295 _3360_ _3439_ _0527_ sky130_fd_sc_hd__o21a_1
X_4346_ VGND VPWR _0050_ _1191_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4277_ VPWR VGND VGND VPWR net69 _1124_ _0844_ sky130_fd_sc_hd__nand2_4
X_7065_ VPWR VGND VPWR VGND _2165_ _3283_ _3334_ _3378_ sky130_fd_sc_hd__or3_1
X_6016_ VGND VPWR VPWR VGND _2574_ i_tinyqv.cpu.instr_data\[2\]\[12\] _2562_ _1712_
+ sky130_fd_sc_hd__mux2_1
X_7967_ i_tinyqv.cpu.i_core.i_registers.rd\[0\] clknet_leaf_5_clk _0104_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6918_ VGND VPWR VPWR VGND _0909_ _0854_ _0956_ _3270_ sky130_fd_sc_hd__or3_2
Xclkbuf_leaf_34_clk VGND VPWR clknet_3_7__leaf_clk clknet_leaf_34_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_7898_ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[21\] clknet_leaf_5_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[21\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6849_ VGND VPWR VPWR VGND _3220_ _3219_ _2991_ _2546_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_508 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_8519_ i_tinyqv.cpu.i_core.i_instrret.register\[25\] clknet_leaf_48_clk i_tinyqv.cpu.i_core.i_instrret.reg_buf\[25\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_490 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_25_clk VGND VPWR clknet_3_6__leaf_clk clknet_leaf_25_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_0_28_538 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_36_560 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xrebuffer3 VPWR VGND VPWR VGND net322 _1412_ sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_11_449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4200_ VPWR VGND _1047_ _1042_ _1040_ VPWR VGND sky130_fd_sc_hd__and2_1
X_5180_ VPWR VGND VGND VPWR _1936_ i_tinyqv.cpu.i_core.multiplier.accum\[11\] _1934_
+ sky130_fd_sc_hd__or2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.i_regbuf\[23\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[23\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[27\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_79_Left_160 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4131_ VPWR VGND VPWR VGND _0978_ i_tinyqv.mem.instr_active sky130_fd_sc_hd__inv_2
X_4062_ VPWR VGND VGND VPWR _0908_ _0909_ _0907_ sky130_fd_sc_hd__nand2_4
Xwire25 VGND VPWR net25 _0671_ VPWR VGND sky130_fd_sc_hd__buf_1
X_7821_ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[8\] clknet_leaf_49_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[8\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4964_ VGND VPWR _1738_ gpio_out\[6\] _1737_ _1730_ VPWR VGND sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_16_clk VGND VPWR clknet_3_2__leaf_clk clknet_leaf_16_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_7752_ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[3\] clknet_leaf_56_clk _0081_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6703_ VGND VPWR VGND VPWR _3087_ _3079_ _3077_ _3076_ sky130_fd_sc_hd__a21bo_1
X_3915_ VGND VPWR _0767_ _0667_ i_tinyqv.cpu.i_core.i_registers.reg_access\[2\]\[1\]
+ _0670_ VPWR VGND sky130_fd_sc_hd__and3_1
X_7683_ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[30\] clknet_leaf_58_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[30\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4895_ VGND VPWR _0062_ _1691_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6634_ VPWR VGND VGND VPWR _1442_ _3026_ _2306_ sky130_fd_sc_hd__nand2_1
X_3846_ VGND VPWR VPWR VGND i_tinyqv.cpu.debug_instr_valid _0698_ i_tinyqv.cpu.is_branch
+ i_tinyqv.cpu.is_alu_reg sky130_fd_sc_hd__o21ai_4
X_6565_ VGND VPWR VPWR VGND _2972_ i_tinyqv.cpu.data_out\[23\] _2912_ i_tinyqv.cpu.data_out\[31\]
+ sky130_fd_sc_hd__mux2_1
X_3777_ VPWR VGND VPWR VGND net53 net56 i_tinyqv.cpu.i_core.i_registers.rs1\[0\] _0629_
+ net52 sky130_fd_sc_hd__or4b_1
X_8304_ i_tinyqv.mem.q_ctrl.data_ready clknet_leaf_16_clk _0403_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_2
X_5516_ VGND VPWR VPWR VGND i_uart_tx.fsm_state\[1\] _2222_ i_uart_tx.fsm_state\[3\]
+ _2223_ i_uart_tx.fsm_state\[0\] sky130_fd_sc_hd__a31oi_1
X_6496_ VGND VPWR VPWR VGND _2910_ i_spi.end_txn _2909_ i_debug_uart_tx.uart_tx_data\[0\]
+ sky130_fd_sc_hd__mux2_1
X_5447_ VPWR VGND VPWR VGND i_uart_tx.cycle_counter\[8\] i_uart_tx.cycle_counter\[7\]
+ i_uart_tx.cycle_counter\[10\] _2173_ i_uart_tx.cycle_counter\[9\] sky130_fd_sc_hd__or4b_1
X_8235_ i_tinyqv.cpu.i_core.mepc\[6\] clknet_leaf_34_clk _0335_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_8166_ i_tinyqv.cpu.instr_data\[2\]\[15\] clknet_leaf_14_clk _0278_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5378_ _2111_ _2083_ _2110_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_8097_ i_tinyqv.cpu.i_core.interrupt_req\[0\] clknet_leaf_26_clk net2 VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_4329_ _1176_ _0742_ _0708_ net78 _1175_ VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_7117_ _3424_ _3292_ _3337_ _3423_ _3304_ VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_7048_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_cycles.rstn _3361_ _3281_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_313 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_9_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xi_tinyqv.cpu.i_core.i_cycles.i_regbuf\[6\] i_tinyqv.cpu.i_core.i_cycles.reg_buf\[6\]
+ i_tinyqv.cpu.i_core.cycle_count_wide\[6\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_56_611 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_28_313 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_4680_ VPWR VGND VGND VPWR _1444_ _1399_ _1516_ _1515_ sky130_fd_sc_hd__nor3_4
X_6350_ VPWR VGND VGND VPWR _2791_ i_tinyqv.mem.q_ctrl.read_cycles_count\[0\] _2782_
+ sky130_fd_sc_hd__or2_1
X_5301_ VGND VPWR _1752_ _2049_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_6281_ VGND VPWR VPWR VGND _2750_ i_tinyqv.cpu.instr_data_in\[5\] _2744_ _1717_ sky130_fd_sc_hd__mux2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.i_regbuf\[24\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[24\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[28\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_8020_ i_uart_rx.fsm_state\[3\] clknet_leaf_30_clk _0155_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_5232_ VPWR VGND VGND VPWR _1984_ _1986_ _1985_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_5_clk VGND VPWR clknet_3_0__leaf_clk clknet_leaf_5_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_5163_ VPWR VGND VGND VPWR _1920_ _1917_ _1918_ sky130_fd_sc_hd__or2_1
X_4114_ VPWR VGND VGND VPWR _0961_ _0959_ _0960_ sky130_fd_sc_hd__or2_1
X_5094_ _1853_ _1849_ _1847_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_4045_ VPWR VGND _0892_ _0891_ i_tinyqv.cpu.instr_data_start\[8\] VPWR VGND sky130_fd_sc_hd__and2_1
Xclone8 VPWR VGND net324 i_tinyqv.cpu.i_core.i_registers.rs1\[3\] VPWR VGND sky130_fd_sc_hd__buf_2
X_7804_ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[23\] clknet_leaf_0_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[23\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5996_ VGND VPWR VPWR VGND _2564_ i_tinyqv.cpu.instr_data\[2\]\[2\] _2563_ i_tinyqv.cpu.instr_data_in\[2\]
+ sky130_fd_sc_hd__mux2_1
X_4947_ VGND VPWR _1726_ _1727_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_7735_ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[18\] clknet_leaf_59_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[18\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_357 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_46_121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_7666_ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[13\] clknet_leaf_56_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[13\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4878_ VGND VPWR VPWR VGND _1682_ i_tinyqv.cpu.debug_rd\[1\] _1680_ net216 sky130_fd_sc_hd__mux2_1
X_6617_ VGND VPWR _2681_ _3012_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_3829_ VGND VPWR VGND VPWR _0662_ _0681_ i_tinyqv.cpu.i_core.i_registers.rs2\[2\]
+ net37 _0661_ sky130_fd_sc_hd__and4bb_2
X_7597_ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[8\] clknet_leaf_0_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[8\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6548_ VPWR VGND VGND VPWR _2316_ _2952_ _2957_ _2958_ sky130_fd_sc_hd__o21a_1
X_6479_ VGND VPWR _0412_ _2899_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8218_ i_tinyqv.cpu.i_core.multiplier.accum\[1\] clknet_leaf_39_clk _0019_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_8149_ VGND VPWR VGND VPWR i_tinyqv.cpu.data_addr\[24\] _0261_ clknet_leaf_40_clk
+ sky130_fd_sc_hd__dfxtp_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.i_regbuf\[12\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[12\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[16\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.i_regbuf\[9\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[9\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[13\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_625 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_80_477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_53_669 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_21_500 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_21_577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xi_tinyqv.cpu.i_core.i_instrret.i_regbuf\[11\] i_tinyqv.cpu.i_core.i_instrret.reg_buf\[11\]
+ i_tinyqv.cpu.i_core.i_instrret.register\[15\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap1 VGND VPWR net320 _0683_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5850_ VPWR VGND _2469_ _2468_ VPWR VGND sky130_fd_sc_hd__buf_4
X_5781_ VPWR VGND VPWR VGND _2384_ _2403_ i_spi.spi_clk_out _2418_ sky130_fd_sc_hd__or3_1
X_4801_ VGND VPWR VGND VPWR _1635_ _0955_ _1636_ _1023_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_0_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_7520_ VPWR VGND _3750_ _3744_ net92 VPWR VGND sky130_fd_sc_hd__and2_1
X_4732_ VGND VPWR VPWR VGND _1565_ _1567_ _1566_ sky130_fd_sc_hd__xor2_1
X_7451_ VGND VPWR VPWR VGND _3696_ _3695_ _3625_ i_tinyqv.mem.q_ctrl.addr\[16\] sky130_fd_sc_hd__mux2_1
XFILLER_0_56_496 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_43_102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_4663_ VGND VPWR VPWR VGND _1499_ i_tinyqv.cpu.instr_data\[3\]\[9\] _1449_ i_tinyqv.cpu.instr_data\[1\]\[9\]
+ sky130_fd_sc_hd__mux2_1
X_6402_ VGND VPWR i_tinyqv.cpu.data_addr\[24\] i_tinyqv.mem.q_ctrl.last_ram_b_sel
+ _2839_ i_tinyqv.cpu.data_addr\[23\] _2734_ VPWR VGND sky130_fd_sc_hd__and4b_1
X_7382_ VPWR VGND VGND VPWR net93 _3624_ _2733_ _3638_ sky130_fd_sc_hd__o21a_1
X_4594_ VPWR VGND VPWR VGND _1422_ i_tinyqv.cpu.instr_write_offset\[2\] _1429_ _1430_
+ sky130_fd_sc_hd__a21o_1
X_6333_ VGND VPWR VPWR VGND _2778_ _1717_ _2772_ net287 sky130_fd_sc_hd__mux2_1
XFILLER_0_12_533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_6264_ VGND VPWR VPWR VGND _1016_ _1531_ _2681_ _2739_ sky130_fd_sc_hd__or3b_1
X_8003_ i_uart_rx.cycle_counter\[7\] clknet_leaf_30_clk _0138_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_5215_ VPWR VGND VGND VPWR _1970_ _1967_ _1968_ sky130_fd_sc_hd__or2_1
X_6195_ VPWR VGND _2679_ _2678_ _1536_ VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_43_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5146_ VGND VPWR _1902_ _1903_ _1878_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_5077_ VGND VPWR _1811_ _1808_ _1837_ _1810_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_4028_ VGND VPWR VPWR VGND _0876_ gpio_out\[4\] gpio_out_sel\[4\] _0875_ sky130_fd_sc_hd__mux2_1
X_5979_ VGND VPWR _0260_ _2551_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7718_ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[1\] clknet_leaf_56_clk _0031_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_603 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7649_ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[28\] clknet_leaf_57_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[28\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.i_regbuf\[24\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[24\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[28\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_190 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.i_regbuf\[13\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[13\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[17\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_48 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_41_617 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold209 net238 i_debug_uart_tx.uart_tx_data\[4\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5000_ VGND VPWR VPWR VGND _1764_ _1440_ _1763_ i_tinyqv.cpu.data_continue sky130_fd_sc_hd__mux2_1
X_6951_ VGND VPWR _3278_ _0612_ _2079_ _0724_ VPWR VGND sky130_fd_sc_hd__and3_1
X_5902_ VGND VPWR VPWR VGND _2499_ _2498_ _2399_ i_spi.data\[7\] sky130_fd_sc_hd__mux2_1
X_6882_ VPWR VGND VPWR VGND _1556_ i_tinyqv.cpu.load_started _1759_ _3246_ sky130_fd_sc_hd__a21o_1
XFILLER_0_64_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.i_regbuf\[4\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[4\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[8\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5833_ VPWR VGND VPWR VGND net230 _2456_ _2457_ _0944_ _2442_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_48_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_29_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_8552_ i_tinyqv.cpu.i_core.i_cycles.register\[25\] clknet_leaf_3_clk i_tinyqv.cpu.i_core.i_cycles.reg_buf\[25\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5764_ VGND VPWR _2404_ net239 _2405_ _2394_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_7503_ VPWR VGND _3739_ _2071_ net121 VPWR VGND sky130_fd_sc_hd__and2_1
X_5695_ VPWR VGND _2351_ _2337_ i_debug_uart_tx.data_to_send\[6\] VPWR VGND sky130_fd_sc_hd__and2_1
X_8483_ i_tinyqv.mem.q_ctrl.addr\[9\] clknet_leaf_32_clk _0581_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_4715_ VPWR VGND VPWR VGND _1551_ _1550_ _1517_ sky130_fd_sc_hd__or2_2
XFILLER_0_17_658 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_7434_ VPWR VGND _3681_ _3676_ i_tinyqv.cpu.instr_data_start\[14\] VPWR VGND sky130_fd_sc_hd__and2_1
X_4646_ VPWR VGND VGND VPWR _1482_ _1481_ _1476_ sky130_fd_sc_hd__or2_1
X_7365_ VGND VPWR _3623_ _1528_ _2079_ _2995_ VPWR VGND sky130_fd_sc_hd__and3_1
X_4577_ VGND VPWR VPWR VGND _1413_ i_tinyqv.cpu.instr_data\[2\]\[0\] net36 i_tinyqv.cpu.instr_data\[0\]\[0\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_691 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6316_ VGND VPWR _0380_ _2768_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7296_ VPWR VGND VPWR VGND _2131_ _3569_ _2142_ _2129_ _3570_ sky130_fd_sc_hd__or4_1
X_6247_ VGND VPWR _2725_ _1813_ _1060_ _2696_ VPWR VGND sky130_fd_sc_hd__and3_1
X_6178_ VGND VPWR VPWR VGND _2670_ i_tinyqv.cpu.i_core.mepc\[16\] _2667_ i_tinyqv.cpu.i_core.mepc\[12\]
+ sky130_fd_sc_hd__mux2_1
X_5129_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.multiplier.accum\[9\] _1887_ _1886_
+ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_24_Left_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_67_514 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_67_569 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_33_Left_114 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_42_Left_123 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold81 net110 i_tinyqv.cpu.data_out\[31\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 net121 i_tinyqv.cpu.i_core.cycle_count\[1\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 net99 i_tinyqv.cpu.i_core.is_double_fault_r VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_51_Left_132 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5480_ VPWR VGND VPWR VGND _2198_ i_debug_uart_tx.resetn sky130_fd_sc_hd__inv_2
X_4500_ VGND VPWR VGND VPWR _1339_ _1206_ _0887_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_14_639 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XANTENNA_1 _0865_ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_4431_ VPWR VGND VGND VPWR _1080_ _1274_ _1273_ sky130_fd_sc_hd__nand2_1
X_4362_ VPWR VGND VGND VPWR _1205_ _0890_ _1204_ sky130_fd_sc_hd__or2_1
X_7150_ VGND VPWR VPWR VGND _1487_ _2125_ _1468_ _3454_ sky130_fd_sc_hd__or3_2
XPHY_EDGE_ROW_60_Left_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4293_ VGND VPWR VPWR VGND _1140_ _1139_ i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt\[1\]
+ _1138_ sky130_fd_sc_hd__mux2_1
X_6101_ VGND VPWR _0315_ _2618_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7081_ VPWR VGND VGND VPWR _3292_ _3349_ _3305_ _3392_ sky130_fd_sc_hd__o21a_1
X_6032_ VGND VPWR VPWR VGND _2582_ i_tinyqv.cpu.instr_data\[1\]\[6\] _2463_ i_tinyqv.cpu.instr_data_in\[6\]
+ sky130_fd_sc_hd__mux2_1
X_7983_ i_uart_tx.cycle_counter\[2\] clknet_leaf_32_clk _0118_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
Xrebuffer46 VGND VPWR net75 net74 VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xrebuffer35 VGND VPWR net64 _0740_ VPWR VGND sky130_fd_sc_hd__buf_1
Xrebuffer24 VGND VPWR net53 i_tinyqv.cpu.i_core.i_registers.rs1\[1\] VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xrebuffer13 VGND VPWR net42 net41 VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6934_ VPWR VGND _3274_ _3273_ VPWR VGND sky130_fd_sc_hd__buf_2
Xrebuffer57 VGND VPWR net86 _0799_ VPWR VGND sky130_fd_sc_hd__buf_1
X_6865_ VGND VPWR _3233_ _3234_ _3232_ VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_569 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_5816_ VPWR VGND VPWR VGND _2443_ _0916_ _2441_ _2444_ sky130_fd_sc_hd__a21oi_1
X_6796_ VPWR VGND VPWR VGND _3164_ _3039_ _3172_ _2306_ _0915_ _3171_ sky130_fd_sc_hd__a221o_1
X_5747_ VGND VPWR _2390_ _2384_ _2181_ _2389_ VPWR VGND sky130_fd_sc_hd__and3_1
X_8535_ i_tinyqv.cpu.i_core.cycle_count_wide\[4\] clknet_leaf_50_clk i_tinyqv.cpu.i_core.i_cycles.reg_buf\[8\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_561 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_8466_ i_tinyqv.cpu.i_core.i_registers.rs2\[1\] clknet_leaf_5_clk _0564_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_32_403 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5678_ VPWR VGND VPWR VGND _2339_ _0989_ sky130_fd_sc_hd__inv_2
X_7417_ VPWR VGND _3667_ _3661_ i_tinyqv.cpu.instr_data_start\[11\] VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_32_436 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_8397_ i_tinyqv.cpu.data_out\[22\] clknet_leaf_20_clk _0495_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.i_regbuf\[27\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[15\].genblk1.genblk1.genblk1.reg_buf\[27\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[15\]\[31\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4629_ VPWR VGND VPWR VGND _1462_ _1461_ _1464_ _1465_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_683 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_7348_ VPWR VGND VGND VPWR i_tinyqv.cpu.additional_mem_ops\[1\] i_tinyqv.cpu.additional_mem_ops\[0\]
+ _3611_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7279_ VPWR VGND VGND VPWR _3337_ _3556_ _3289_ sky130_fd_sc_hd__nor2_2
XFILLER_0_79_193 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_63_561 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_78_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_4980_ VPWR VGND VPWR VGND _1741_ net238 _1747_ _0012_ sky130_fd_sc_hd__a21o_1
XFILLER_0_53_78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_3931_ VGND VPWR VGND VPWR _0781_ _0747_ _0783_ _0782_ sky130_fd_sc_hd__a21oi_2
X_6650_ VPWR VGND VPWR VGND _3038_ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[12\]
+ sky130_fd_sc_hd__inv_2
X_3862_ VPWR VGND VGND VPWR _0714_ _0713_ _0712_ _0710_ _0709_ sky130_fd_sc_hd__nor4_1
X_5601_ VPWR VGND VGND VPWR _1228_ _2283_ _2282_ sky130_fd_sc_hd__nand2_1
X_6581_ VGND VPWR VPWR VGND _2983_ _2982_ _2562_ i_tinyqv.cpu.instr_data_in\[1\] sky130_fd_sc_hd__mux2_1
X_5532_ VGND VPWR VGND VPWR i_uart_rx.cycle_counter\[2\] i_uart_rx.cycle_counter\[4\]
+ i_uart_rx.cycle_counter\[5\] i_uart_rx.cycle_counter\[3\] _2235_ sky130_fd_sc_hd__and4bb_1
X_8320_ i_tinyqv.cpu.instr_data_in\[8\] clknet_leaf_16_clk _0419_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_3793_ VGND VPWR VGND VPWR i_tinyqv.cpu.i_core.i_registers.rs1\[1\] i_tinyqv.cpu.i_core.i_registers.rs1\[3\]
+ i_tinyqv.cpu.i_core.i_registers.rs1\[2\] i_tinyqv.cpu.i_core.i_registers.rs1\[0\]
+ _0645_ sky130_fd_sc_hd__and4bb_1
X_8251_ debug_register_data clknet_leaf_19_clk _0351_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_5463_ VGND VPWR VGND VPWR _0110_ net98 _2169_ _2186_ _2182_ sky130_fd_sc_hd__o211a_1
X_8182_ i_tinyqv.cpu.i_core.i_shift.a\[1\] clknet_leaf_41_clk _0294_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
X_4414_ VPWR VGND VGND VPWR _1257_ _1255_ _1256_ sky130_fd_sc_hd__or2_1
X_5394_ VGND VPWR _1476_ _2124_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_7202_ VPWR VGND VGND VPWR _2126_ _3351_ _3298_ _3498_ sky130_fd_sc_hd__o21a_1
X_7133_ VGND VPWR VGND VPWR _3439_ _3434_ _3437_ _3364_ _3438_ sky130_fd_sc_hd__a211o_1
X_4345_ VGND VPWR VPWR VGND _1191_ i_tinyqv.cpu.debug_rd\[0\] _1190_ i_tinyqv.cpu.i_core.i_registers.reg_access\[15\]\[0\]
+ sky130_fd_sc_hd__mux2_1
X_4276_ VPWR VGND VGND VPWR _1030_ _1123_ _1122_ sky130_fd_sc_hd__nand2_1
X_7064_ _3300_ _3299_ _3377_ _2121_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_6015_ VGND VPWR _0274_ _2573_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_620 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_7966_ i_tinyqv.cpu.i_core.mstatus_mte clknet_leaf_37_clk _0103_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_6917_ VGND VPWR VPWR VGND _0480_ _3269_ _3265_ _1619_ _3266_ net273 sky130_fd_sc_hd__a32o_1
X_7897_ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[20\] clknet_leaf_48_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[20\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6848_ VGND VPWR _3218_ _3219_ _3217_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_6779_ VPWR VGND _3156_ _3146_ _3148_ VPWR VGND sky130_fd_sc_hd__and2_1
X_8518_ i_tinyqv.cpu.i_core.i_instrret.register\[24\] clknet_leaf_50_clk i_tinyqv.cpu.i_core.i_instrret.reg_buf\[24\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.i_regbuf\[28\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[28\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_8449_ i_tinyqv.cpu.imm\[27\] clknet_leaf_8_clk _0547_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.i_regbuf\[31\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[31\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[3\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xrebuffer4 VGND VPWR net33 _1397_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.i_regbuf\[27\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[27\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[31\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_cycles.i_regbuf\[25\] i_tinyqv.cpu.i_core.i_cycles.reg_buf\[25\]
+ i_tinyqv.cpu.i_core.i_cycles.register\[29\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4130_ VPWR VGND _0977_ _0872_ i_tinyqv.mem.q_ctrl.data_ready VPWR VGND sky130_fd_sc_hd__and2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.i_regbuf\[16\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[16\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[20\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4061_ VGND VPWR VPWR VGND _0838_ _0908_ sky130_fd_sc_hd__clkinv_4
X_7820_ i_tinyqv.cpu.i_core.i_registers.reg_access\[6\]\[3\] clknet_leaf_52_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[7\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4963_ VPWR VGND _1737_ _1728_ VPWR VGND sky130_fd_sc_hd__buf_2
X_7751_ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[2\] clknet_leaf_1_clk _0080_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6702_ VPWR VGND VGND VPWR _3084_ _3086_ _3085_ sky130_fd_sc_hd__nand2_1
X_7682_ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[29\] clknet_leaf_57_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[29\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_3914_ VGND VPWR VGND VPWR _0766_ net61 _0764_ i_tinyqv.cpu.i_core.i_registers.reg_access\[14\]\[1\]
+ _0765_ sky130_fd_sc_hd__a211o_1
XFILLER_0_74_645 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_6633_ VGND VPWR VPWR VGND _0440_ _3025_ _3024_ _3005_ _3009_ net95 sky130_fd_sc_hd__a32o_1
X_4894_ VGND VPWR VPWR VGND _1691_ _1184_ _1690_ i_tinyqv.cpu.i_core.i_registers.reg_access\[5\]\[0\]
+ sky130_fd_sc_hd__mux2_1
X_3845_ VGND VPWR _0696_ _0688_ _0697_ _0693_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_13_70 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_6564_ VGND VPWR _0425_ _2971_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_3776_ VGND VPWR net324 _0624_ _0628_ _0627_ _0625_ VPWR VGND sky130_fd_sc_hd__and4b_1
X_8303_ i_tinyqv.mem.q_ctrl.fsm_state\[2\] clknet_leaf_15_clk _0402_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5515_ VPWR VGND VPWR VGND _2222_ i_uart_tx.fsm_state\[2\] sky130_fd_sc_hd__inv_2
X_6495_ VPWR VGND _2909_ _2908_ VPWR VGND sky130_fd_sc_hd__buf_2
X_5446_ VPWR VGND VPWR VGND i_uart_tx.cycle_counter\[4\] i_uart_tx.cycle_counter\[6\]
+ _2172_ i_uart_tx.cycle_counter\[5\] i_uart_tx.cycle_counter\[3\] sky130_fd_sc_hd__or4bb_1
X_8234_ i_tinyqv.cpu.i_core.mepc\[5\] clknet_leaf_40_clk _0334_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_8165_ i_tinyqv.cpu.instr_data\[2\]\[14\] clknet_leaf_12_clk _0277_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5377_ VGND VPWR VPWR VGND _2110_ i_tinyqv.cpu.i_core.mstatus_mpie _2109_ _2104_
+ sky130_fd_sc_hd__mux2_1
X_8096_ gpio_out\[7\] clknet_leaf_17_clk _0007_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4328_ net69 _0656_ _1175_ _1030_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_7116_ VPWR VGND VPWR VGND _3423_ _3415_ sky130_fd_sc_hd__inv_2
X_4259_ VGND VPWR VPWR VGND _1106_ i_tinyqv.cpu.i_core.i_shift.a\[11\] _1028_ i_tinyqv.cpu.i_core.i_shift.a\[20\]
+ sky130_fd_sc_hd__mux2_1
X_7047_ VGND VPWR _3359_ _3360_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_7949_ i_tinyqv.cpu.i_core.mcause\[0\] clknet_leaf_37_clk _0087_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_394 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_34_58 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_51_350 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_3_425 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5300_ VPWR VGND _0085_ _1604_ i_tinyqv.cpu.i_core.cycle\[0\] _1753_ _2048_ VGND
+ VPWR sky130_fd_sc_hd__a31o_1
X_6280_ VGND VPWR _0363_ _2749_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5231_ VPWR VGND VGND VPWR _1985_ i_tinyqv.cpu.i_core.multiplier.accum\[13\] _1983_
+ sky130_fd_sc_hd__or2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.i_regbuf\[17\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[17\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[21\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5162_ VPWR VGND VGND VPWR _1917_ _1919_ _1918_ sky130_fd_sc_hd__nand2_1
X_4113_ VPWR VGND VPWR VGND i_tinyqv.cpu.data_addr\[26\] i_tinyqv.cpu.data_addr\[25\]
+ i_tinyqv.cpu.data_addr\[0\] _0960_ i_tinyqv.cpu.data_addr\[27\] sky130_fd_sc_hd__or4b_1
X_5093_ VPWR VGND VGND VPWR _1851_ _1852_ _0021_ sky130_fd_sc_hd__nor2_1
X_4044_ VGND VPWR _0891_ _0883_ i_tinyqv.cpu.instr_data_start\[7\] _0890_ VPWR VGND
+ sky130_fd_sc_hd__and3_1
X_7803_ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[22\] clknet_leaf_57_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[22\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5995_ VPWR VGND _2563_ _2562_ VPWR VGND sky130_fd_sc_hd__buf_4
X_7734_ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[17\] clknet_leaf_55_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[17\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4946_ VPWR VGND _1726_ _1725_ _1001_ VPWR VGND sky130_fd_sc_hd__and2_1
X_7665_ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[12\] clknet_leaf_0_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[12\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.i_regbuf\[20\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[20\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[24\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4877_ VGND VPWR _0070_ _1681_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6616_ VGND VPWR VPWR VGND _3011_ _2988_ _3010_ _1406_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_230 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_15_520 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7596_ i_tinyqv.cpu.i_core.i_registers.reg_access\[13\]\[3\] clknet_leaf_1_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[7\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_3828_ VGND VPWR VGND VPWR net37 _0680_ i_tinyqv.cpu.i_core.i_registers.rs2\[3\]
+ net38 i_tinyqv.cpu.i_core.i_registers.rs2\[2\] sky130_fd_sc_hd__and4bb_2
X_6547_ VGND VPWR VGND VPWR _2957_ _2953_ _2955_ _2914_ _2956_ sky130_fd_sc_hd__a211o_1
XFILLER_0_6_285 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_15_564 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_3759_ VGND VPWR _0607_ _0611_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_6478_ VGND VPWR VPWR VGND _2899_ net133 _2897_ net11 sky130_fd_sc_hd__mux2_1
X_5429_ VGND VPWR VPWR VGND _2158_ i_tinyqv.cpu.i_core.i_registers.rd\[1\] _2153_
+ _2157_ sky130_fd_sc_hd__mux2_1
X_8217_ i_tinyqv.cpu.i_core.multiplier.accum\[0\] clknet_leaf_39_clk _0016_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_589 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_8148_ VGND VPWR VGND VPWR i_tinyqv.cpu.data_addr\[23\] _0260_ clknet_leaf_35_clk
+ sky130_fd_sc_hd__dfxtp_4
X_8079_ debug_rd_r\[3\] clknet_leaf_53_clk net32 VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_648 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_53_637 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_40_309 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_21_534 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xmax_cap2 VGND VPWR net321 _0634_ VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_0_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_206 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_4800_ _1635_ _1620_ _1624_ _1630_ _1634_ VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_0_61_23 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5780_ VPWR VGND VPWR VGND _1725_ _1000_ _2386_ _2417_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_528 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_29_656 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4731_ VPWR VGND VGND VPWR _0701_ _1566_ _0820_ sky130_fd_sc_hd__nand2_1
X_7450_ VGND VPWR VPWR VGND _3695_ _3694_ _3004_ net147 sky130_fd_sc_hd__mux2_1
XFILLER_0_4_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_4662_ VGND VPWR VPWR VGND _1498_ _1497_ _1409_ _1496_ sky130_fd_sc_hd__mux2_1
X_6401_ VPWR VGND VPWR VGND i_tinyqv.cpu.data_addr\[24\] _2838_ i_tinyqv.cpu.data_addr\[23\]
+ _2681_ sky130_fd_sc_hd__or3b_2
XFILLER_0_9_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_7381_ VGND VPWR VGND VPWR _3637_ net299 _2682_ _3004_ _3636_ sky130_fd_sc_hd__o211a_1
X_4593_ VGND VPWR _1428_ _1429_ i_tinyqv.cpu.instr_write_offset\[3\] VPWR VGND sky130_fd_sc_hd__xnor2_1
X_6332_ VGND VPWR _0387_ _2777_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_191 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_12_556 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_6263_ VGND VPWR _0357_ _2738_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8002_ i_uart_rx.cycle_counter\[6\] clknet_leaf_30_clk _0137_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_5214_ VPWR VGND VGND VPWR _1967_ _1969_ _1968_ sky130_fd_sc_hd__nand2_1
X_6194_ VPWR VGND VGND VPWR _1551_ _1541_ _2678_ sky130_fd_sc_hd__nor2_1
X_5145_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_shift.a\[8\] _1902_ _1880_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5076_ VGND VPWR VPWR VGND _1834_ _1836_ _1835_ sky130_fd_sc_hd__xor2_1
X_4027_ VGND VPWR VPWR VGND debug_register_data debug_rd_r\[2\] i_spi.spi_select _0875_
+ sky130_fd_sc_hd__mux2_2
XFILLER_0_79_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.i_regbuf\[21\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[21\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[25\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5978_ VGND VPWR VPWR VGND _2551_ _2550_ _2501_ i_tinyqv.cpu.data_addr\[23\] sky130_fd_sc_hd__mux2_1
X_4929_ VGND VPWR VGND VPWR i_tinyqv.mem.q_ctrl.fsm_state\[1\] _1714_ _1707_ sky130_fd_sc_hd__or2b_1
X_7717_ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[0\] clknet_leaf_1_clk _0030_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_453 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_7648_ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[27\] clknet_leaf_46_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[27\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.i_regbuf\[7\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[7\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[11\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7579_ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[22\] clknet_leaf_55_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[22\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.i_regbuf\[10\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[10\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[14\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.i_regbuf\[17\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[17\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[21\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.i_regbuf\[5\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[5\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[9\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_442 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_53_434 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_41_607 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_6950_ VPWR VGND VGND VPWR _2066_ _0974_ _0505_ sky130_fd_sc_hd__nor2_1
X_5901_ VGND VPWR VPWR VGND _2498_ i_spi.data\[6\] _2386_ i_debug_uart_tx.uart_tx_data\[7\]
+ sky130_fd_sc_hd__mux2_1
X_6881_ VGND VPWR VGND VPWR _0468_ _1762_ _3245_ net258 _2067_ sky130_fd_sc_hd__a211o_1
X_5832_ VPWR VGND VPWR VGND _2088_ _1312_ _2434_ _2456_ sky130_fd_sc_hd__a21o_1
X_5763_ _2392_ _2404_ i_spi.spi_clk_out _2403_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_8551_ i_tinyqv.cpu.i_core.i_cycles.register\[24\] clknet_leaf_51_clk i_tinyqv.cpu.i_core.i_cycles.reg_buf\[24\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4714_ VPWR VGND VGND VPWR _1550_ _1480_ _1546_ sky130_fd_sc_hd__or2_1
X_7502_ _0596_ net248 i_tinyqv.cpu.i_core.cycle_count\[0\] _0744_ _3738_ VPWR VGND
+ VGND VPWR sky130_fd_sc_hd__o31a_1
X_5694_ VGND VPWR VGND VPWR _0177_ i_debug_uart_tx.uart_tx_data\[4\] _2330_ _2350_
+ _2299_ sky130_fd_sc_hd__o211a_1
X_8482_ i_tinyqv.mem.q_ctrl.addr\[8\] clknet_leaf_33_clk _0580_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_136 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7433_ VPWR VGND VGND VPWR _3680_ i_tinyqv.cpu.instr_data_start\[14\] _3676_ sky130_fd_sc_hd__or2_1
X_4645_ VPWR VGND VPWR VGND _1470_ _1416_ _1472_ _1481_ sky130_fd_sc_hd__a21o_1
X_4576_ VGND VPWR VPWR VGND _1339_ _1410_ _1412_ _1411_ sky130_fd_sc_hd__o21a_4
X_7364_ VPWR VGND _0574_ _2066_ _3622_ _1410_ _3619_ _3618_ VPWR VGND sky130_fd_sc_hd__a311oi_1
X_6315_ VGND VPWR VPWR VGND _2768_ _1717_ _2762_ i_tinyqv.mem.data_from_read\[21\]
+ sky130_fd_sc_hd__mux2_1
X_7295_ VPWR VGND VGND VPWR _1483_ _2122_ _3569_ sky130_fd_sc_hd__nor2_1
X_6246_ VGND VPWR _2724_ _0354_ _2714_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_6177_ VGND VPWR _0340_ _2669_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5128_ VGND VPWR VPWR VGND _1884_ _1886_ _1885_ sky130_fd_sc_hd__xor2_1
X_5059_ VGND VPWR VPWR VGND _1817_ _1820_ _1819_ sky130_fd_sc_hd__xor2_1
XFILLER_0_47_261 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_35_445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold60 net89 i_tinyqv.mem.q_ctrl.addr\[6\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 net111 i_tinyqv.cpu.data_addr\[14\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 net100 i_tinyqv.cpu.instr_data\[3\]\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 net122 i_tinyqv.mem.q_ctrl.addr\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.i_regbuf\[21\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[21\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[25\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_261 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XANTENNA_2 _0991_ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_4430_ VGND VPWR VPWR VGND _1273_ _1095_ _1149_ _1073_ sky130_fd_sc_hd__mux2_1
X_4361_ VPWR VGND VGND VPWR i_tinyqv.cpu.instr_data_start\[5\] _0889_ _1204_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_6100_ VGND VPWR VPWR VGND _2618_ i_tinyqv.cpu.i_core.i_shift.a\[22\] _2595_ i_tinyqv.cpu.i_core.i_shift.a\[26\]
+ sky130_fd_sc_hd__mux2_1
X_4292_ VGND VPWR VPWR VGND _1139_ _1105_ _1050_ _1102_ sky130_fd_sc_hd__mux2_1
X_7080_ VGND VPWR VPWR VGND _3391_ _3390_ _3319_ _1501_ sky130_fd_sc_hd__mux2_1
X_6031_ VGND VPWR _0282_ _2581_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7982_ i_uart_tx.cycle_counter\[1\] clknet_leaf_31_clk _0117_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
Xrebuffer25 VGND VPWR net54 _0642_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xrebuffer36 VGND VPWR net65 _0740_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xrebuffer14 VGND VPWR net43 _0652_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6933_ VPWR VGND VGND VPWR _0854_ _3263_ _3273_ sky130_fd_sc_hd__nor2_1
Xrebuffer47 VGND VPWR net76 _0793_ VPWR VGND sky130_fd_sc_hd__buf_1
Xrebuffer58 VGND VPWR net87 i_tinyqv.cpu.i_core.i_registers.rs1\[0\] VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6864_ VGND VPWR i_tinyqv.cpu.imm\[23\] _3233_ i_tinyqv.cpu.instr_data_start\[23\]
+ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_5815_ VGND VPWR VGND VPWR i_tinyqv.cpu.i_core.last_interrupt_req\[0\] _2443_ i_tinyqv.cpu.i_core.interrupt_req\[0\]
+ sky130_fd_sc_hd__or2b_1
X_6795_ VGND VPWR VGND VPWR _3171_ _3040_ _3169_ _3170_ _3047_ sky130_fd_sc_hd__o211a_1
X_5746_ VGND VPWR _2385_ _2389_ i_spi.clock_count\[1\] VPWR VGND sky130_fd_sc_hd__xnor2_1
X_8534_ i_tinyqv.cpu.i_core.cycle_count\[3\] clknet_leaf_50_clk i_tinyqv.cpu.i_core.i_cycles.reg_buf\[7\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5677_ VPWR VGND _2338_ _2337_ i_debug_uart_tx.data_to_send\[1\] VPWR VGND sky130_fd_sc_hd__and2_1
X_8465_ i_tinyqv.cpu.i_core.i_registers.rs2\[0\] clknet_leaf_52_clk _0563_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_0_44_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_7416_ VPWR VGND VGND VPWR _3666_ i_tinyqv.cpu.instr_data_start\[11\] _3661_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_448 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_4628_ VGND VPWR VGND VPWR _1464_ i_tinyqv.cpu.instr_data\[0\]\[4\] _1414_ _1409_
+ _1463_ sky130_fd_sc_hd__o211a_1
X_8396_ i_tinyqv.cpu.data_out\[21\] clknet_leaf_20_clk _0494_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_7347_ VPWR VGND _3610_ _3563_ _2124_ _3291_ _3609_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_4559_ VGND VPWR VGND VPWR _1392_ _1394_ _1395_ i_tinyqv.cpu.i_core.is_interrupt
+ sky130_fd_sc_hd__a21oi_2
X_7278_ VPWR VGND VGND VPWR _3293_ _3322_ _3555_ sky130_fd_sc_hd__nor2_1
X_6229_ VPWR VGND VGND VPWR _2709_ _2706_ _2707_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_710 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_2_309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_53_35 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_3930_ VPWR VGND VGND VPWR _0763_ _0780_ _0782_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_356 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_3861_ VPWR VGND VPWR VGND _0678_ i_tinyqv.cpu.i_core.i_registers.reg_access\[11\]\[0\]
+ _0664_ _0713_ i_tinyqv.cpu.i_core.i_registers.reg_access\[7\]\[0\] sky130_fd_sc_hd__a22o_1
X_5600_ VPWR VGND VGND VPWR _0997_ _2282_ _1558_ sky130_fd_sc_hd__nand2_1
X_6580_ VPWR VGND VGND VPWR _2982_ _1400_ i_tinyqv.cpu.instr_data\[2\]\[1\] sky130_fd_sc_hd__or2_1
X_3792_ VPWR VGND _0644_ _0643_ i_tinyqv.cpu.i_core.i_registers.reg_access\[14\]\[3\]
+ VPWR VGND sky130_fd_sc_hd__and2_1
X_5531_ VPWR VGND VGND VPWR net165 _2234_ _0130_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_551 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_6_659 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_8250_ i_tinyqv.cpu.i_core.load_top_bit clknet_leaf_22_clk _0350_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_14_437 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_78_32 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5462_ VPWR VGND VGND VPWR _2186_ _2179_ _2185_ sky130_fd_sc_hd__or2_1
X_7201_ VPWR VGND _3497_ _3496_ _3290_ VPWR VGND sky130_fd_sc_hd__and2_1
X_8181_ i_tinyqv.cpu.i_core.i_shift.a\[0\] clknet_leaf_42_clk _0293_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
X_4413_ VGND VPWR VGND VPWR _0782_ _1256_ _0781_ sky130_fd_sc_hd__or2b_1
X_5393_ VGND VPWR _1481_ _2123_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_4344_ i_tinyqv.cpu.i_core.i_registers.rd\[0\] _1190_ i_tinyqv.cpu.i_core.i_registers.rd\[1\]
+ _1189_ VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_7132_ VGND VPWR _3361_ _3438_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_676 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7063_ VPWR VGND _3376_ _3375_ _3364_ VPWR VGND sky130_fd_sc_hd__and2_1
X_6014_ VGND VPWR VPWR VGND _2573_ i_tinyqv.cpu.instr_data\[2\]\[11\] _2563_ _2322_
+ sky130_fd_sc_hd__mux2_1
X_4275_ VPWR VGND _1122_ _1119_ _1079_ _1046_ _1121_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_7965_ i_tinyqv.cpu.i_core.mstatus_mie clknet_leaf_37_clk _0102_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_6916_ VPWR VGND VGND VPWR _3260_ _3269_ net50 sky130_fd_sc_hd__nor2_2
X_7896_ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[19\] clknet_leaf_48_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[19\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6847_ VGND VPWR _3207_ _3209_ _3218_ _3208_ VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_6778_ VPWR VGND VGND VPWR _3153_ _3155_ _3154_ sky130_fd_sc_hd__nand2_1
X_5729_ _2375_ i_debug_uart_tx.fsm_state\[0\] i_debug_uart_tx.fsm_state\[2\] i_debug_uart_tx.fsm_state\[1\]
+ _2333_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
X_8517_ i_tinyqv.cpu.i_core.i_instrret.register\[23\] clknet_leaf_46_clk i_tinyqv.cpu.i_core.i_instrret.reg_buf\[23\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_510 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_5_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_8448_ i_tinyqv.cpu.imm\[26\] clknet_leaf_7_clk _0546_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_8379_ i_debug_uart_tx.uart_tx_data\[4\] clknet_leaf_19_clk _0477_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.i_regbuf\[24\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[24\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[28\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_49 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xrebuffer5 VGND VPWR net34 net36 VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xi_tinyqv.cpu.i_core.i_cycles.i_regbuf\[18\] i_tinyqv.cpu.i_core.i_cycles.reg_buf\[18\]
+ i_tinyqv.cpu.i_core.i_cycles.register\[22\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4060_ _0907_ _0614_ VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xwire16 VPWR VGND net16 _0808_ VPWR VGND sky130_fd_sc_hd__buf_4
X_4962_ VPWR VGND VPWR VGND _1727_ i_debug_uart_tx.uart_tx_data\[5\] _1736_ _0005_
+ sky130_fd_sc_hd__a21o_1
X_7750_ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[1\] clknet_leaf_55_clk _0079_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6701_ VPWR VGND VGND VPWR _3085_ i_tinyqv.cpu.instr_data_start\[8\] i_tinyqv.cpu.i_core.imm_lo\[8\]
+ sky130_fd_sc_hd__or2_1
X_7681_ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[28\] clknet_leaf_59_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[28\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_3913_ VPWR VGND VPWR VGND _0680_ i_tinyqv.cpu.i_core.i_registers.reg_access\[15\]\[1\]
+ _0677_ _0765_ i_tinyqv.cpu.i_core.i_registers.reg_access\[9\]\[1\] sky130_fd_sc_hd__a22o_1
X_4893_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.i_registers.rd\[3\] _1188_ _1647_
+ i_tinyqv.cpu.i_core.i_registers.rd\[2\] _1690_ sky130_fd_sc_hd__and4b_2
X_6632_ VPWR VGND VGND VPWR _3025_ i_tinyqv.cpu.data_addr\[3\] _3012_ sky130_fd_sc_hd__or2_1
X_3844_ VGND VPWR VGND VPWR _0696_ _0689_ _0695_ i_tinyqv.cpu.imm\[19\] _0611_ sky130_fd_sc_hd__a211o_1
X_6563_ VGND VPWR VPWR VGND _2971_ _1720_ _2925_ _2970_ sky130_fd_sc_hd__mux2_1
X_3775_ VPWR VGND _0627_ i_tinyqv.cpu.i_core.i_registers.rs1\[0\] VPWR VGND sky130_fd_sc_hd__buf_4
X_8302_ i_tinyqv.mem.q_ctrl.fsm_state\[1\] clknet_leaf_15_clk _0401_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
X_5514_ VGND VPWR _1728_ _2221_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_6494_ VPWR VGND _2908_ _2907_ _2906_ VPWR VGND sky130_fd_sc_hd__and2_1
X_5445_ VPWR VGND VGND VPWR net206 _2171_ i_uart_tx.cycle_counter\[0\] sky130_fd_sc_hd__nand2_1
X_8233_ i_tinyqv.cpu.i_core.mepc\[4\] clknet_leaf_35_clk _0333_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_8164_ i_tinyqv.cpu.instr_data\[2\]\[13\] clknet_leaf_12_clk _0276_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_7115_ VGND VPWR _0525_ _3422_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5376_ VPWR VGND VGND VPWR _2109_ _2057_ _2108_ _2107_ _1348_ _0939_ sky130_fd_sc_hd__o41a_1
X_8095_ gpio_out\[6\] clknet_leaf_18_clk _0006_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4327_ VGND VPWR VGND VPWR _1173_ _1171_ _0745_ _1174_ sky130_fd_sc_hd__o21ba_1
X_4258_ VGND VPWR VPWR VGND _1105_ i_tinyqv.cpu.i_core.i_shift.a\[10\] _1028_ i_tinyqv.cpu.i_core.i_shift.a\[21\]
+ sky130_fd_sc_hd__mux2_1
X_7046_ VPWR VGND _3359_ _3358_ VPWR VGND sky130_fd_sc_hd__buf_2
X_4189_ VPWR VGND _1036_ _1027_ VPWR VGND sky130_fd_sc_hd__buf_4
X_7948_ i_tinyqv.cpu.i_core.cycle\[1\] clknet_leaf_51_clk _0086_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_7879_ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[2\] clknet_leaf_5_clk _0064_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_189 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold190 net219 i_uart_tx.cycle_counter\[3\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.i_regbuf\[25\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[25\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[29\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_16_Right_16 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_25_Right_25 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5230_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.multiplier.accum\[13\] _1984_ _1983_
+ sky130_fd_sc_hd__nand2_1
X_5161_ VGND VPWR _1893_ _1890_ _1918_ _1892_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_4112_ VPWR VGND VPWR VGND i_tinyqv.cpu.data_addr\[1\] i_tinyqv.cpu.data_addr\[6\]
+ i_tinyqv.cpu.data_addr\[7\] i_tinyqv.cpu.data_addr\[24\] _0959_ sky130_fd_sc_hd__or4_1
X_5092_ VPWR VGND VGND VPWR _1850_ _1827_ _1830_ _1852_ sky130_fd_sc_hd__nor3_1
X_4043_ VPWR VGND _0890_ _0889_ i_tinyqv.cpu.instr_data_start\[5\] VPWR VGND sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_34_Right_34 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5994_ VGND VPWR _2561_ _2562_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_7802_ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[21\] clknet_leaf_1_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[21\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4945_ VGND VPWR _1557_ _1725_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_7733_ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[16\] clknet_leaf_59_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[16\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7664_ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[11\] clknet_leaf_45_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[11\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4876_ VGND VPWR VPWR VGND _1681_ i_tinyqv.cpu.debug_rd\[0\] _1680_ i_tinyqv.cpu.i_core.i_registers.reg_access\[7\]\[0\]
+ sky130_fd_sc_hd__mux2_1
X_6615_ VGND VPWR i_tinyqv.cpu.was_early_branch _3010_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.i_regbuf\[13\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[13\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[17\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3827_ VPWR VGND VPWR VGND _0678_ i_tinyqv.cpu.i_core.i_registers.reg_access\[15\]\[3\]
+ _0677_ _0679_ i_tinyqv.cpu.i_core.i_registers.reg_access\[7\]\[3\] sky130_fd_sc_hd__a22o_1
X_7595_ i_tinyqv.cpu.i_core.i_registers.reg_access\[13\]\[2\] clknet_leaf_2_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[6\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_43_Right_43 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6546_ VPWR VGND VGND VPWR _2956_ _1713_ _2916_ sky130_fd_sc_hd__nand2_2
X_3758_ VPWR VGND VGND VPWR _0609_ _0610_ _0607_ sky130_fd_sc_hd__nor2_2
XFILLER_0_40_80 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_15_587 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6477_ VGND VPWR _0411_ _2898_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5428_ _2157_ _2147_ _1641_ _1647_ _2156_ VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_8216_ i_tinyqv.cpu.i_core.i_shift.b\[3\] clknet_leaf_39_clk _0328_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5359_ VGND VPWR _1395_ _2094_ _2095_ _0754_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_8147_ i_tinyqv.cpu.data_addr\[22\] clknet_leaf_34_clk _0259_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_8078_ debug_rd_r\[2\] clknet_leaf_51_clk i_tinyqv.cpu.debug_rd\[2\] VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_52_Right_52 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_7029_ _0517_ _3340_ _3343_ _3344_ _2061_ VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
XPHY_EDGE_ROW_61_Right_61 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_70_Right_70 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_29_668 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4730_ VPWR VGND VGND VPWR _0817_ _1565_ _1324_ sky130_fd_sc_hd__nand2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.i_regbuf\[8\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[8\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[12\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4661_ VGND VPWR VPWR VGND _1497_ i_tinyqv.cpu.instr_data\[2\]\[10\] _1449_ i_tinyqv.cpu.instr_data\[0\]\[10\]
+ sky130_fd_sc_hd__mux2_1
X_6400_ VPWR VGND VGND VPWR _2794_ _2836_ _2837_ sky130_fd_sc_hd__nor2_1
X_7380_ VPWR VGND VPWR VGND _3632_ _3056_ _3636_ _3633_ _3635_ _2877_ sky130_fd_sc_hd__a221o_1
X_6331_ VGND VPWR VPWR VGND _2777_ _1712_ _2772_ net276 sky130_fd_sc_hd__mux2_1
X_4592_ VPWR VGND VGND VPWR _0653_ _1428_ _0888_ sky130_fd_sc_hd__nand2_1
X_6262_ VGND VPWR _2738_ _2733_ _2181_ _2737_ VPWR VGND sky130_fd_sc_hd__and3_1
X_8001_ i_uart_rx.cycle_counter\[5\] clknet_leaf_30_clk _0136_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_5213_ VGND VPWR _1941_ _1938_ _1968_ _1940_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_6193_ VGND VPWR _0348_ _2677_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5144_ VPWR VGND VGND VPWR _1884_ _1901_ _1885_ sky130_fd_sc_hd__nand2_1
X_5075_ VPWR VGND VGND VPWR _1054_ _1835_ _1167_ sky130_fd_sc_hd__nand2_1
X_4026_ VPWR VGND uo_out[0] _0874_ VPWR VGND sky130_fd_sc_hd__buf_4
X_5977_ VGND VPWR VPWR VGND _2550_ i_tinyqv.cpu.i_core.mepc\[23\] _2504_ i_tinyqv.cpu.i_core.i_shift.a\[27\]
+ sky130_fd_sc_hd__mux2_1
X_4928_ VGND VPWR i_tinyqv.mem.q_ctrl.is_writing _1713_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_7716_ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[31\] clknet_leaf_59_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[31\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.i_regbuf\[14\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[6\].genblk1.genblk1.genblk1.reg_buf\[14\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[6\]\[18\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7647_ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[26\] clknet_leaf_46_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[26\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4859_ VGND VPWR VPWR VGND _1671_ i_tinyqv.cpu.debug_rd\[1\] _1669_ net254 sky130_fd_sc_hd__mux2_1
X_7578_ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[21\] clknet_leaf_58_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[21\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_0__f_clk VGND VPWR VGND VPWR clknet_0_clk clknet_3_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_6529_ VGND VPWR VPWR VGND _2941_ _2940_ _2920_ net12 sky130_fd_sc_hd__mux2_1
XFILLER_0_43_682 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_8_Left_89 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.i_regbuf\[7\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[7\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[11\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_421 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.i_regbuf\[5\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[5\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[9\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_321 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5900_ VGND VPWR _0235_ _2497_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6880_ VPWR VGND VGND VPWR i_tinyqv.cpu.data_write_n\[1\] _1556_ _3243_ _3245_ sky130_fd_sc_hd__o21a_1
X_5831_ VPWR VGND VPWR VGND _2455_ _2454_ _2083_ _0209_ sky130_fd_sc_hd__a21oi_1
X_5762_ VPWR VGND VPWR VGND i_spi.bits_remaining\[2\] _2402_ i_spi.bits_remaining\[3\]
+ _2403_ sky130_fd_sc_hd__or3_1
XFILLER_0_8_326 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_8550_ i_tinyqv.cpu.i_core.i_cycles.register\[23\] clknet_leaf_50_clk i_tinyqv.cpu.i_core.i_cycles.reg_buf\[23\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4713_ VPWR VGND VPWR VGND _1545_ _1384_ _1549_ _1548_ net8 sky130_fd_sc_hd__a211oi_2
X_7501_ VPWR VGND VGND VPWR _2066_ _2071_ _3738_ sky130_fd_sc_hd__nor2_1
X_5693_ VGND VPWR VGND VPWR _2350_ _2336_ _2341_ i_debug_uart_tx.data_to_send\[4\]
+ _2349_ sky130_fd_sc_hd__a211o_1
X_8481_ i_tinyqv.mem.q_ctrl.addr\[7\] clknet_leaf_32_clk _0579_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_7432_ VPWR VGND VPWR VGND net187 _3007_ _0585_ _3009_ net304 _3679_ sky130_fd_sc_hd__a221o_1
X_4644_ VPWR VGND VGND VPWR _1444_ _1399_ _1480_ _1479_ sky130_fd_sc_hd__nor3_4
X_4575_ VPWR VGND VPWR VGND _1411_ i_tinyqv.cpu.debug_instr_valid i_tinyqv.cpu.pc\[2\]
+ sky130_fd_sc_hd__or2_2
X_7363_ VGND VPWR VPWR VGND _3622_ _3619_ _3618_ _2993_ _3621_ sky130_fd_sc_hd__o2bb2a_1
X_6314_ VGND VPWR _0379_ _2767_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7294_ VGND VPWR _0558_ _3568_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6245_ _2724_ _2722_ _2723_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_6176_ VGND VPWR VPWR VGND _2669_ i_tinyqv.cpu.i_core.mepc\[15\] _2667_ i_tinyqv.cpu.i_core.mepc\[11\]
+ sky130_fd_sc_hd__mux2_1
X_5127_ VGND VPWR _1855_ _1857_ _1885_ _1831_ VPWR VGND sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_2_Right_2 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5058_ VPWR VGND VPWR VGND _1796_ i_tinyqv.cpu.i_core.multiplier.accum\[5\] _1818_
+ _1819_ sky130_fd_sc_hd__a21o_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.i_regbuf\[4\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[4\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[8\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4009_ VPWR VGND _0860_ _0851_ _0849_ i_tinyqv.cpu.i_core.load_done _0859_ VGND VPWR
+ sky130_fd_sc_hd__a31o_1
Xhold83 net112 i_tinyqv.cpu.data_out\[21\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 net101 i_tinyqv.cpu.i_core.i_registers.reg_access\[12\]\[3\] VPWR VGND VGND
+ VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 VGND VPWR net90 i_tinyqv.cpu.i_core.i_instrret.data\[3\] VPWR VGND sky130_fd_sc_hd__buf_1
Xhold94 net123 i_tinyqv.cpu.i_core.mcause\[3\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_55_clk VGND VPWR clknet_3_1__leaf_clk clknet_leaf_55_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.i_regbuf\[14\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[1\].genblk1.genblk1.genblk1.reg_buf\[14\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[1\]\[18\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_424 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_13_107 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_41_438 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XANTENNA_3 _1054_ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_4360_ VPWR VGND VPWR VGND _1203_ _1202_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4291_ VGND VPWR VPWR VGND _1138_ _1101_ _1050_ _1137_ sky130_fd_sc_hd__mux2_1
X_6030_ VGND VPWR VPWR VGND _2581_ i_tinyqv.cpu.instr_data\[1\]\[5\] _2463_ i_tinyqv.cpu.instr_data_in\[5\]
+ sky130_fd_sc_hd__mux2_1
X_7981_ i_uart_tx.cycle_counter\[0\] clknet_leaf_32_clk _0116_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
Xrebuffer26 VGND VPWR net55 _0649_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xrebuffer15 VGND VPWR net44 net20 VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6932_ VPWR VGND VPWR VGND _3272_ _3253_ _3269_ _0492_ net143 sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_46_clk VGND VPWR clknet_3_4__leaf_clk clknet_leaf_46_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xrebuffer59 VGND VPWR net88 _0649_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xrebuffer48 VGND VPWR net77 _0720_ VPWR VGND sky130_fd_sc_hd__buf_1
Xrebuffer37 VGND VPWR _0762_ net66 VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_6863_ VGND VPWR _3224_ _3226_ _3232_ _3225_ VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_112 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5814_ VPWR VGND VGND VPWR _1312_ _2102_ _2442_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_6794_ VPWR VGND VGND VPWR _1390_ _3170_ _2536_ sky130_fd_sc_hd__nand2_1
X_5745_ VGND VPWR _0190_ _2388_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8533_ i_tinyqv.cpu.i_core.cycle_count\[2\] clknet_leaf_51_clk i_tinyqv.cpu.i_core.i_cycles.reg_buf\[6\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5676_ VGND VPWR _2337_ _2333_ _0988_ _2335_ VPWR VGND sky130_fd_sc_hd__and3_1
X_8464_ i_tinyqv.cpu.i_core.i_registers.rs1\[3\] clknet_leaf_51_clk _0562_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_7415_ VPWR VGND VPWR VGND net89 _3007_ _0582_ _3009_ net317 _3665_ sky130_fd_sc_hd__a221o_1
X_4627_ VPWR VGND VGND VPWR _1463_ i_tinyqv.cpu.instr_data\[2\]\[4\] _1422_ sky130_fd_sc_hd__or2_1
X_8395_ i_tinyqv.cpu.data_out\[20\] clknet_leaf_19_clk _0493_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_7346_ VPWR VGND VPWR VGND _1514_ _2143_ _3609_ _3351_ _2155_ _2149_ sky130_fd_sc_hd__a221o_1
X_4558_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.imm_lo\[8\] i_tinyqv.cpu.i_core.imm_lo\[9\]
+ _1394_ sky130_fd_sc_hd__nor2_1
X_4489_ VGND VPWR VPWR VGND _1328_ _0828_ _1178_ _0827_ _1327_ sky130_fd_sc_hd__o2bb2a_1
X_7277_ VPWR VGND VPWR VGND _3554_ _3553_ sky130_fd_sc_hd__inv_2
X_6228_ VPWR VGND _2708_ _2707_ _2706_ VPWR VGND sky130_fd_sc_hd__and2_1
X_6159_ VGND VPWR VPWR VGND _2660_ i_tinyqv.cpu.i_core.mepc\[7\] _2656_ i_tinyqv.cpu.i_core.mepc\[3\]
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_37_clk VGND VPWR clknet_3_4__leaf_clk clknet_leaf_37_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_0_63_585 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_28_clk VGND VPWR clknet_3_6__leaf_clk clknet_leaf_28_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_0_58_379 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_3860_ _0712_ _0711_ i_tinyqv.cpu.counter\[4\] _0620_ _0670_ VGND VPWR VPWR VGND
+ sky130_fd_sc_hd__and4_1
X_3791_ VGND VPWR net51 i_tinyqv.cpu.i_core.i_registers.rs1\[0\] _0643_ net30 net70
+ VPWR VGND sky130_fd_sc_hd__and4b_1
X_5530_ VGND VPWR _2225_ _2233_ i_uart_tx.fsm_state\[1\] _2234_ _2198_ i_uart_tx.fsm_state\[3\]
+ VPWR VGND sky130_fd_sc_hd__a41o_1
X_5461_ VGND VPWR VPWR VGND _2185_ i_uart_tx.data_to_send\[3\] _2177_ i_uart_tx.data_to_send\[2\]
+ sky130_fd_sc_hd__mux2_1
X_7200_ VPWR VGND VPWR VGND i_tinyqv.cpu.instr_data\[0\]\[1\] _3487_ _3496_ _3488_
+ i_tinyqv.cpu.instr_data\[1\]\[1\] _3495_ sky130_fd_sc_hd__a221o_1
X_4412_ VPWR VGND VPWR VGND _0745_ _0743_ _0746_ _1255_ sky130_fd_sc_hd__a21oi_1
X_8180_ i_tinyqv.cpu.instr_data\[1\]\[15\] clknet_leaf_11_clk _0292_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5392_ VPWR VGND VPWR VGND _2122_ _1469_ _1486_ sky130_fd_sc_hd__or2_2
X_4343_ VGND VPWR _1189_ i_tinyqv.cpu.i_core.i_registers.rd\[3\] i_tinyqv.cpu.i_core.i_registers.rd\[2\]
+ _1188_ VPWR VGND sky130_fd_sc_hd__and3_1
X_7131_ VPWR VGND VPWR VGND _1514_ _3352_ _3437_ _3435_ _2155_ _3436_ sky130_fd_sc_hd__a221o_1
X_4274_ _1121_ _1046_ _1120_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_7062_ VGND VPWR VPWR VGND _3375_ _3374_ _3319_ _1467_ _3320_ _1510_ sky130_fd_sc_hd__a32o_1
X_6013_ VGND VPWR _0273_ _2572_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_19_clk VGND VPWR clknet_3_3__leaf_clk clknet_leaf_19_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_7964_ i_tinyqv.cpu.i_core.mstatus_mpie clknet_leaf_38_clk _0101_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_633 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6915_ VGND VPWR VPWR VGND _0479_ _3268_ _3265_ _1619_ _3266_ net234 sky130_fd_sc_hd__a32o_1
XFILLER_0_11_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_7895_ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[18\] clknet_leaf_3_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[18\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6846_ VPWR VGND VGND VPWR _3215_ _3217_ _3216_ sky130_fd_sc_hd__nand2_1
X_6777_ VPWR VGND VGND VPWR _3154_ _0881_ i_tinyqv.cpu.imm\[15\] sky130_fd_sc_hd__or2_1
X_5728_ VGND VPWR _0187_ _2374_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8516_ i_tinyqv.cpu.i_core.i_instrret.register\[22\] clknet_leaf_48_clk i_tinyqv.cpu.i_core.i_instrret.reg_buf\[22\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_3989_ VPWR VGND _0840_ _0839_ VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_0_60_522 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_8447_ i_tinyqv.cpu.imm\[25\] clknet_leaf_9_clk _0545_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5659_ VGND VPWR VPWR VGND _2324_ _1712_ _2308_ i_tinyqv.cpu.instr_data\[3\]\[12\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_693 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_8378_ i_debug_uart_tx.uart_tx_data\[3\] clknet_leaf_26_clk _0476_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_2
X_7329_ VPWR VGND VGND VPWR _3595_ _3596_ _3597_ sky130_fd_sc_hd__nor2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.i_regbuf\[28\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[28\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.i_regbuf\[17\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[17\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[21\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xrebuffer6 VGND VPWR net35 net36 VPWR VGND sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_39_Left_120 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xi_tinyqv.cpu.i_core.i_instrret.i_regbuf\[27\] i_tinyqv.cpu.i_core.i_instrret.reg_buf\[27\]
+ i_tinyqv.cpu.i_core.i_instrret.register\[31\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xwire17 VGND VPWR net17 _2241_ VPWR VGND sky130_fd_sc_hd__buf_1
Xwire28 VPWR VGND net28 _0972_ VPWR VGND sky130_fd_sc_hd__buf_2
X_4961_ VGND VPWR _1736_ gpio_out\[5\] _1729_ _1730_ VPWR VGND sky130_fd_sc_hd__and3_1
X_6700_ VPWR VGND VGND VPWR i_tinyqv.cpu.instr_data_start\[8\] _3084_ i_tinyqv.cpu.i_core.imm_lo\[8\]
+ sky130_fd_sc_hd__nand2_1
X_7680_ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[27\] clknet_leaf_46_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[27\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4892_ VGND VPWR _0069_ _1689_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_3912_ VPWR VGND VPWR VGND _0674_ i_tinyqv.cpu.i_core.i_registers.reg_access\[8\]\[1\]
+ _0671_ _0764_ i_tinyqv.cpu.i_core.i_registers.reg_access\[12\]\[1\] sky130_fd_sc_hd__a22o_1
X_6631_ VPWR VGND VPWR VGND _3016_ _3018_ _3024_ _3023_ _3017_ _2878_ sky130_fd_sc_hd__a221o_1
X_3843_ VPWR VGND VPWR VGND i_tinyqv.cpu.imm\[23\] _0619_ _0695_ _0690_ i_tinyqv.cpu.imm\[27\]
+ _0694_ sky130_fd_sc_hd__a221o_1
X_8301_ i_tinyqv.mem.q_ctrl.fsm_state\[0\] clknet_leaf_15_clk _0400_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_6562_ VPWR VGND VGND VPWR _2320_ _2952_ _2969_ _2970_ sky130_fd_sc_hd__o21a_1
X_3774_ VPWR VGND _0626_ i_tinyqv.cpu.i_core.i_registers.rs1\[3\] VPWR VGND sky130_fd_sc_hd__buf_6
X_5513_ VPWR VGND VPWR VGND _2218_ net102 _2220_ _0126_ sky130_fd_sc_hd__a21oi_1
X_6493_ VPWR VGND VGND VPWR _2907_ _0868_ i_tinyqv.mem.q_ctrl.data_req sky130_fd_sc_hd__or2_1
XFILLER_0_42_533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5444_ VGND VPWR i_uart_tx.fsm_state\[1\] i_uart_tx.fsm_state\[3\] _2170_ i_uart_tx.fsm_state\[2\]
+ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_8232_ i_tinyqv.cpu.i_core.mepc\[3\] clknet_leaf_35_clk _0332_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_8_clk VGND VPWR clknet_3_3__leaf_clk clknet_leaf_8_clk VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_8163_ i_tinyqv.cpu.instr_data\[2\]\[12\] clknet_leaf_11_clk _0275_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_7114_ VGND VPWR VPWR VGND _3422_ _3421_ _3396_ i_tinyqv.cpu.i_core.imm_lo\[5\] sky130_fd_sc_hd__mux2_1
X_5375_ VGND VPWR _0652_ _0920_ _2108_ _0844_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_8094_ gpio_out\[5\] clknet_leaf_17_clk _0005_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4326_ VPWR VGND VGND VPWR _1173_ _0843_ _0919_ sky130_fd_sc_hd__nand2_2
X_4257_ VGND VPWR VPWR VGND _1104_ _1102_ _1103_ _1101_ sky130_fd_sc_hd__mux2_1
X_7045_ VPWR VGND VGND VPWR _1400_ _3295_ _3358_ sky130_fd_sc_hd__nor2_1
X_4188_ VPWR VGND VPWR VGND _1025_ i_tinyqv.cpu.i_core.cmp _1034_ _1035_ sky130_fd_sc_hd__a21o_1
X_7947_ i_tinyqv.cpu.i_core.cycle\[0\] clknet_leaf_51_clk _0085_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_2
X_7878_ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[1\] clknet_leaf_53_clk _0063_
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6829_ VPWR VGND VGND VPWR _2987_ _1601_ _3202_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold180 net209 i_tinyqv.cpu.is_system VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 net220 i_spi.read_latency VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.i_regbuf\[29\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[29\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[1\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.i_regbuf\[18\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[8\].genblk1.genblk1.genblk1.reg_buf\[18\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[8\]\[22\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_522 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xi_tinyqv.cpu.i_core.i_cycles.i_regbuf\[30\] i_tinyqv.cpu.i_core.i_cycles.reg_buf\[30\]
+ i_tinyqv.cpu.i_core.i_cycles.register\[2\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5160_ VGND VPWR VPWR VGND _1915_ _1917_ _1916_ sky130_fd_sc_hd__xor2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.i_regbuf\[21\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[21\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[13\]\[25\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4111_ VPWR VGND VPWR VGND i_tinyqv.mem.data_from_read\[16\] _0689_ _0958_ _0748_
+ i_tinyqv.mem.data_from_read\[20\] _0957_ sky130_fd_sc_hd__a221o_1
X_5091_ VPWR VGND VGND VPWR _1830_ _1827_ _1850_ _1851_ sky130_fd_sc_hd__o21a_1
X_4042_ VGND VPWR _0889_ _0884_ i_tinyqv.cpu.instr_data_start\[4\] _0888_ VPWR VGND
+ sky130_fd_sc_hd__and3_1
X_5993_ VGND VPWR VPWR VGND _2460_ i_tinyqv.cpu.instr_write_offset\[2\] _1406_ _2561_
+ sky130_fd_sc_hd__or3b_1
X_7801_ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[20\] clknet_leaf_3_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[20\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4944_ VGND VPWR _1724_ uio_oe[5] VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_7732_ i_tinyqv.cpu.i_core.i_registers.registers\[9\]\[15\] clknet_leaf_53_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[9\].genblk1.genblk1.genblk1.reg_buf\[15\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_7663_ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[10\] clknet_leaf_58_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[10\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_4875_ VPWR VGND VGND VPWR _1679_ _1680_ _1188_ i_tinyqv.cpu.i_core.i_registers.rd\[3\]
+ sky130_fd_sc_hd__nor3b_2
X_6614_ VGND VPWR VPWR VGND _0437_ _3005_ _2878_ net300 _3009_ net122 sky130_fd_sc_hd__a32o_1
X_7594_ i_tinyqv.cpu.i_core.i_registers.reg_access\[13\]\[1\] clknet_leaf_53_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[13\].genblk1.genblk1.genblk1.reg_buf\[5\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_3826_ VPWR VGND VGND VPWR _0661_ i_tinyqv.cpu.i_core.i_registers.rs2\[2\] net37
+ net38 _0678_ sky130_fd_sc_hd__and4b_2
X_6545_ VGND VPWR VGND VPWR _2955_ i_tinyqv.cpu.data_out\[12\] _2912_ _2929_ _2954_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_190 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_3757_ VGND VPWR VGND VPWR i_tinyqv.cpu.counter\[3\] _0609_ _0608_ sky130_fd_sc_hd__or2b_1
X_6476_ VGND VPWR VPWR VGND _2898_ i_tinyqv.mem.q_ctrl.spi_in_buffer\[0\] _2897_ net10
+ sky130_fd_sc_hd__mux2_1
X_8215_ i_tinyqv.cpu.i_core.i_shift.b\[2\] clknet_leaf_39_clk _0327_ VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_5427_ VPWR VGND VPWR VGND _1514_ _2137_ _2156_ _2141_ _2155_ _2149_ sky130_fd_sc_hd__a221o_1
X_5358_ VGND VPWR VGND VPWR _2094_ net18 _2093_ net66 _2056_ sky130_fd_sc_hd__a211o_1
X_8146_ i_tinyqv.cpu.data_addr\[21\] clknet_leaf_35_clk _0258_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_8077_ debug_rd_r\[1\] clknet_leaf_52_clk i_tinyqv.cpu.debug_rd\[1\] VPWR VGND VPWR
+ VGND sky130_fd_sc_hd__dfxtp_1
X_4309_ VGND VPWR VPWR VGND _1156_ _1155_ _1108_ _1154_ sky130_fd_sc_hd__mux2_1
X_5289_ VPWR VGND VGND VPWR _2039_ _2041_ _2040_ sky130_fd_sc_hd__nand2_1
X_7028_ _2155_ _1466_ _3344_ _3333_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
XFILLER_0_37_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_53_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xi_tinyqv.cpu.i_core.i_cycles.i_regbuf\[4\] i_tinyqv.cpu.i_core.i_cycles.reg_buf\[4\]
+ i_tinyqv.cpu.i_core.cycle_count_wide\[4\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_56_444 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4660_ VGND VPWR VPWR VGND _1496_ i_tinyqv.cpu.instr_data\[3\]\[10\] _1449_ i_tinyqv.cpu.instr_data\[1\]\[10\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_330 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_6330_ VGND VPWR _0386_ _2776_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4591_ VPWR VGND VPWR VGND _1427_ _1420_ _1426_ sky130_fd_sc_hd__or2_2
XFILLER_0_3_213 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_6261_ VGND VPWR VPWR VGND _2737_ _2735_ _0868_ _2736_ sky130_fd_sc_hd__mux2_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.i_regbuf\[22\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[7\].genblk1.genblk1.genblk1.reg_buf\[22\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[7\]\[26\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_8000_ i_uart_rx.cycle_counter\[4\] clknet_leaf_31_clk _0135_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.i_regbuf\[8\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[8\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[12\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5212_ VGND VPWR VPWR VGND _1965_ _1967_ _1966_ sky130_fd_sc_hd__xor2_1
X_6192_ VGND VPWR VPWR VGND _2677_ i_tinyqv.cpu.i_core.mepc\[23\] _2667_ i_tinyqv.cpu.i_core.mepc\[19\]
+ sky130_fd_sc_hd__mux2_1
X_5143_ VGND VPWR VPWR VGND _1899_ _0023_ _1900_ sky130_fd_sc_hd__xor2_1
X_5074_ VPWR VGND VGND VPWR _1832_ _1834_ _1833_ sky130_fd_sc_hd__nand2_1
X_4025_ VGND VPWR VPWR VGND _0874_ gpio_out\[0\] gpio_out_sel\[0\] i_uart_tx.txd_reg
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_35_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5976_ VGND VPWR _0259_ _2549_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_4927_ VGND VPWR i_tinyqv.cpu.instr_data_in\[12\] _1712_ VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_7715_ i_tinyqv.cpu.i_core.i_registers.registers\[10\]\[30\] clknet_leaf_56_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[10\].genblk1.genblk1.genblk1.reg_buf\[30\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_285 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_62_425 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_62_414 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_4858_ VGND VPWR _0078_ _1670_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_7646_ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[25\] clknet_leaf_57_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[25\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_3809_ VPWR VGND _0661_ i_tinyqv.cpu.i_core.i_registers.rs2\[3\] VPWR VGND sky130_fd_sc_hd__buf_2
X_4789_ VGND VPWR VGND VPWR _1624_ _0957_ _1623_ _0971_ _0907_ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_7577_ i_tinyqv.cpu.i_core.i_registers.registers\[14\]\[20\] clknet_leaf_59_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[14\].genblk1.genblk1.genblk1.reg_buf\[20\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_6528_ VGND VPWR VPWR VGND _2940_ i_tinyqv.mem.q_ctrl.spi_in_buffer\[2\] _2918_ i_tinyqv.mem.q_ctrl.spi_in_buffer\[6\]
+ sky130_fd_sc_hd__mux2_1
X_6459_ VPWR VGND VPWR VGND _2792_ i_tinyqv.mem.q_ctrl.spi_flash_select _1708_ _2884_
+ sky130_fd_sc_hd__a21o_1
X_8129_ i_tinyqv.cpu.data_addr\[4\] clknet_leaf_28_clk _0241_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.i_regbuf\[10\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[11\].genblk1.genblk1.genblk1.reg_buf\[10\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[11\]\[14\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.i_regbuf\[7\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[7\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[11\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_76_506 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_5830_ VGND VPWR VPWR VGND net67 _0944_ _2102_ _2455_ sky130_fd_sc_hd__or3b_1
X_5761_ VPWR VGND VGND VPWR _2402_ i_spi.bits_remaining\[1\] i_spi.bits_remaining\[0\]
+ sky130_fd_sc_hd__or2_1
XFILLER_0_8_305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4712_ VPWR VGND VGND VPWR _1384_ _1547_ _1548_ sky130_fd_sc_hd__nor2_1
X_7500_ VGND VPWR _0595_ _3737_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_8480_ i_tinyqv.mem.q_ctrl.addr\[6\] clknet_leaf_33_clk _0578_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_5692_ VPWR VGND _2349_ _2337_ i_debug_uart_tx.data_to_send\[5\] VPWR VGND sky130_fd_sc_hd__and2_1
X_7431_ VGND VPWR VGND VPWR _3679_ net181 _3012_ _3004_ _3678_ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_499 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_4643_ VGND VPWR VGND VPWR _1478_ _1427_ _1467_ _1479_ sky130_fd_sc_hd__o21ba_1
X_4574_ VPWR VGND VPWR VGND _1410_ i_tinyqv.cpu.debug_instr_valid sky130_fd_sc_hd__inv_2
X_7362_ VPWR VGND VGND VPWR _2150_ _3621_ _1515_ sky130_fd_sc_hd__nand2_1
X_6313_ VGND VPWR VPWR VGND _2767_ _1712_ _2762_ net292 sky130_fd_sc_hd__mux2_1
XFILLER_0_12_344 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_7293_ VGND VPWR VPWR VGND _3568_ _3567_ _3395_ i_tinyqv.cpu.i_core.mem_op\[2\] sky130_fd_sc_hd__mux2_1
X_6244_ VPWR VGND VGND VPWR _2704_ _2723_ _2721_ sky130_fd_sc_hd__nand2_1
X_6175_ VGND VPWR _0339_ _2668_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5126_ VGND VPWR VPWR VGND _1882_ _1884_ _1883_ sky130_fd_sc_hd__xor2_1
X_5057_ VPWR VGND _1818_ _1795_ _1793_ VPWR VGND sky130_fd_sc_hd__and2_1
X_4008_ VPWR VGND VPWR VGND _0837_ _0857_ _0858_ _0859_ _0856_ sky130_fd_sc_hd__nand4_1
XFILLER_0_1_71 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_39_219 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_5959_ VGND VPWR VPWR VGND _2538_ i_tinyqv.cpu.i_core.mepc\[17\] _2504_ i_tinyqv.cpu.i_core.i_shift.a\[21\]
+ sky130_fd_sc_hd__mux2_1
X_7629_ i_tinyqv.cpu.i_core.i_registers.registers\[12\]\[8\] clknet_leaf_56_clk i_tinyqv.cpu.i_core.i_registers.genblk1\[12\].genblk1.genblk1.genblk1.reg_buf\[8\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_35_458 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.i_regbuf\[22\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[2\].genblk1.genblk1.genblk1.reg_buf\[22\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[2\]\[26\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xi_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.i_regbuf\[11\]
+ i_tinyqv.cpu.i_core.i_registers.genblk1\[5\].genblk1.genblk1.genblk1.reg_buf\[11\]
+ i_tinyqv.cpu.i_core.i_registers.registers\[5\]\[15\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 net91 i_uart_rx.cycle_counter\[0\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 net102 i_uart_tx.cycle_counter\[10\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 net113 i_tinyqv.cpu.data_out\[23\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 net124 i_tinyqv.cpu.data_out\[27\] VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_244 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Left_101 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XANTENNA_4 _1185_ VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_0_22_675 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4290_ VGND VPWR VPWR VGND _1137_ _1054_ _1036_ i_tinyqv.cpu.i_core.i_shift.a\[24\]
+ sky130_fd_sc_hd__mux2_1
X_7980_ i_uart_tx.data_to_send\[7\] clknet_leaf_28_clk _0115_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
Xrebuffer16 VGND VPWR net45 net44 VPWR VGND sky130_fd_sc_hd__buf_1
Xrebuffer27 VGND VPWR net56 i_tinyqv.cpu.i_core.i_registers.rs1\[3\] VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6931_ VPWR VGND VPWR VGND _3272_ _3253_ _3268_ _0491_ net175 sky130_fd_sc_hd__a22o_1
Xrebuffer49 VGND VPWR net78 net77 VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xrebuffer38 VGND VPWR net67 net66 VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_6862_ VGND VPWR VGND VPWR _0463_ i_tinyqv.cpu.instr_data_start\[22\] _3123_ _3231_
+ _3205_ sky130_fd_sc_hd__o211a_1
X_5813_ VPWR VGND _2441_ _2088_ _1312_ _0613_ _2435_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_6793_ VGND VPWR _3168_ _3169_ _3165_ VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_403 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_8532_ i_tinyqv.cpu.i_core.cycle_count\[1\] clknet_leaf_6_clk i_tinyqv.cpu.i_core.i_cycles.reg_buf\[5\]
+ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_5744_ _2388_ _2385_ _1729_ _2384_ _2387_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
X_5675_ VGND VPWR VGND VPWR _2335_ _0988_ _2336_ _2333_ sky130_fd_sc_hd__nand3_4
X_8463_ i_tinyqv.cpu.i_core.i_registers.rs1\[2\] clknet_leaf_51_clk _0561_ VPWR VGND
+ VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_8394_ i_tinyqv.cpu.data_out\[19\] clknet_leaf_26_clk _0492_ VPWR VGND VPWR VGND
+ sky130_fd_sc_hd__dfxtp_1
X_7414_ VPWR VGND VGND VPWR net298 _2682_ _3664_ _3665_ sky130_fd_sc_hd__o21a_1
X_4626_ VGND VPWR VPWR VGND _1462_ i_tinyqv.cpu.instr_data\[3\]\[4\] _1414_ i_tinyqv.cpu.instr_data\[1\]\[4\]
+ sky130_fd_sc_hd__mux2_1
X_7345_ VPWR VGND VPWR VGND _3608_ _3607_ _2067_ _0569_ sky130_fd_sc_hd__a21oi_1
X_4557_ VPWR VGND VGND VPWR i_tinyqv.cpu.i_core.imm_lo\[8\] i_tinyqv.cpu.i_core.imm_lo\[9\]
+ _1393_ _1392_ sky130_fd_sc_hd__nand3_1
X_4488_ VGND VPWR VGND VPWR _1175_ _0828_ _1177_ _1327_ sky130_fd_sc_hd__o21ba_1
X_7276_ VPWR VGND VGND VPWR _1473_ _1493_ _3553_ sky130_fd_sc_hd__nor2_1
X_6227_ VGND VPWR _2038_ _2036_ _2707_ _2037_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_6158_ VGND VPWR _0331_ _2659_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_5109_ VGND VPWR VPWR VGND _1866_ _1868_ _1867_ sky130_fd_sc_hd__xor2_1
X_6089_ VGND VPWR _0309_ _2612_ VPWR VGND sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_11_Left_92 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_3790_ VGND VPWR VGND VPWR _0624_ _0642_ net324 _0627_ _0625_ sky130_fd_sc_hd__and4bb_2
X_5460_ VGND VPWR VGND VPWR _0109_ net97 _2169_ _2184_ _2182_ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_417 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_4411_ VGND VPWR VGND VPWR _1254_ _0779_ _0763_ _1175_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_1_322 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_5391_ VPWR VGND _2121_ _2120_ VPWR VGND sky130_fd_sc_hd__buf_2
X_4342_ VGND VPWR VGND VPWR _1186_ _1187_ _1188_ _0877_ sky130_fd_sc_hd__a21oi_4
X_7130_ VPWR VGND VGND VPWR _1507_ _3346_ _3347_ _3334_ _3436_ sky130_fd_sc_hd__o22ai_1
X_4273_ VPWR VGND VGND VPWR i_tinyqv.cpu.alu_op\[3\] _1120_ i_tinyqv.cpu.i_core.i_shift.a\[31\]
+ sky130_fd_sc_hd__nand2_1
X_7061_ VPWR VGND VGND VPWR _3368_ i_tinyqv.cpu.instr_data\[1\]\[4\] _3366_ i_tinyqv.cpu.instr_data\[0\]\[4\]
+ _3374_ _3373_ sky130_fd_sc_hd__o221a_2
X_6012_ VGND VPWR VPWR VGND _2572_ i_tinyqv.cpu.instr_data\[2\]\[10\] _2563_ _2320_
+ sky130_fd_sc_hd__mux2_1
.ends

